`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09.12.2020 11:50:51
// Design Name: 
// Module Name: filterbanks
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module filterbanks(
    input clk,
    input rst,
    input [31:0] powspectr,
    input tvalid_powspectr,
    
    output reg [31:0] feat_filterbanks,
    output reg tvalid_feat_filterbanks
    );
    
    reg [31:0] powspectr_temp;
    reg tvalid_powspectr_temp = 1'b0;
    
    reg [0:25] tvalid_reg_fb;
    reg [31:0] reg_fb_1;
    reg [31:0] reg_fb_2;
    reg [31:0] reg_fb_3;
    reg [31:0] reg_fb_4;
    reg [31:0] reg_fb_5;
    reg [31:0] reg_fb_6;
    reg [31:0] reg_fb_7;
    reg [31:0] reg_fb_8;
    reg [31:0] reg_fb_9;
    reg [31:0] reg_fb_10;
    reg [31:0] reg_fb_11;
    reg [31:0] reg_fb_12;
    reg [31:0] reg_fb_13;
    reg [31:0] reg_fb_14;
    reg [31:0] reg_fb_15;
    reg [31:0] reg_fb_16;
    reg [31:0] reg_fb_17;
    reg [31:0] reg_fb_18;
    reg [31:0] reg_fb_19;
    reg [31:0] reg_fb_20;
    reg [31:0] reg_fb_21;
    reg [31:0] reg_fb_22;
    reg [31:0] reg_fb_23;
    reg [31:0] reg_fb_24;
    reg [31:0] reg_fb_25;
    reg [31:0] reg_fb_26;
    
    reg [11:0] ind = 0;
    
    wire [31:0] filter_banks_1 [0:256];
    wire [31:0] filter_banks_2 [0:256];
    wire [31:0] filter_banks_3 [0:256];
    wire [31:0] filter_banks_4 [0:256];
    wire [31:0] filter_banks_5 [0:256];
    wire [31:0] filter_banks_6 [0:256];
    wire [31:0] filter_banks_7 [0:256];
    wire [31:0] filter_banks_8 [0:256];
    wire [31:0] filter_banks_9 [0:256];
    wire [31:0] filter_banks_10 [0:256];
    wire [31:0] filter_banks_11 [0:256];
    wire [31:0] filter_banks_12 [0:256];
    wire [31:0] filter_banks_13 [0:256];
    wire [31:0] filter_banks_14 [0:256];
    wire [31:0] filter_banks_15 [0:256];
    wire [31:0] filter_banks_16 [0:256];
    wire [31:0] filter_banks_17 [0:256];
    wire [31:0] filter_banks_18 [0:256];
    wire [31:0] filter_banks_19 [0:256];
    wire [31:0] filter_banks_20 [0:256];
    wire [31:0] filter_banks_21 [0:256];
    wire [31:0] filter_banks_22 [0:256];
    wire [31:0] filter_banks_23 [0:256];
    wire [31:0] filter_banks_24 [0:256];
    wire [31:0] filter_banks_25 [0:256];
    wire [31:0] filter_banks_26 [0:256];
    
    
    wire [0:25] tvalid_res_mult_fb;
    wire [31:0] res_mult_fb_1;
    wire [31:0] res_mult_fb_2;
    wire [31:0] res_mult_fb_3;
    wire [31:0] res_mult_fb_4;
    wire [31:0] res_mult_fb_5;
    wire [31:0] res_mult_fb_6;
    wire [31:0] res_mult_fb_7;
    wire [31:0] res_mult_fb_8;
    wire [31:0] res_mult_fb_9;
    wire [31:0] res_mult_fb_10;
    wire [31:0] res_mult_fb_11;
    wire [31:0] res_mult_fb_12;
    wire [31:0] res_mult_fb_13;
    wire [31:0] res_mult_fb_14;
    wire [31:0] res_mult_fb_15;
    wire [31:0] res_mult_fb_16;
    wire [31:0] res_mult_fb_17;
    wire [31:0] res_mult_fb_18;
    wire [31:0] res_mult_fb_19;
    wire [31:0] res_mult_fb_20;
    wire [31:0] res_mult_fb_21;
    wire [31:0] res_mult_fb_22;
    wire [31:0] res_mult_fb_23;
    wire [31:0] res_mult_fb_24;
    wire [31:0] res_mult_fb_25;
    wire [31:0] res_mult_fb_26;
    
    wire [0:25] tvalid_res_add_fb;
    wire [31:0] res_add_fb_1;
    wire [31:0] res_add_fb_2;
    wire [31:0] res_add_fb_3;
    wire [31:0] res_add_fb_4;
    wire [31:0] res_add_fb_5;
    wire [31:0] res_add_fb_6;
    wire [31:0] res_add_fb_7;
    wire [31:0] res_add_fb_8;
    wire [31:0] res_add_fb_9;
    wire [31:0] res_add_fb_10;
    wire [31:0] res_add_fb_11;
    wire [31:0] res_add_fb_12;
    wire [31:0] res_add_fb_13;
    wire [31:0] res_add_fb_14;
    wire [31:0] res_add_fb_15;
    wire [31:0] res_add_fb_16;
    wire [31:0] res_add_fb_17;
    wire [31:0] res_add_fb_18;
    wire [31:0] res_add_fb_19;
    wire [31:0] res_add_fb_20;
    wire [31:0] res_add_fb_21;
    wire [31:0] res_add_fb_22;
    wire [31:0] res_add_fb_23;
    wire [31:0] res_add_fb_24;
    wire [31:0] res_add_fb_25;
    wire [31:0] res_add_fb_26; 
    
    reg [0:25] tvalid_out_acc;
    reg [31:0] out_acc_1;
    reg [31:0] out_acc_2;
    reg [31:0] out_acc_3;
    reg [31:0] out_acc_4;
    reg [31:0] out_acc_5;
    reg [31:0] out_acc_6;
    reg [31:0] out_acc_7;
    reg [31:0] out_acc_8;
    reg [31:0] out_acc_9;
    reg [31:0] out_acc_10;
    reg [31:0] out_acc_11;
    reg [31:0] out_acc_12;
    reg [31:0] out_acc_13;
    reg [31:0] out_acc_14;
    reg [31:0] out_acc_15;
    reg [31:0] out_acc_16;
    reg [31:0] out_acc_17;
    reg [31:0] out_acc_18;
    reg [31:0] out_acc_19;
    reg [31:0] out_acc_20;
    reg [31:0] out_acc_21;
    reg [31:0] out_acc_22;
    reg [31:0] out_acc_23;
    reg [31:0] out_acc_24;
    reg [31:0] out_acc_25;
    reg [31:0] out_acc_26;
    
    reg [31:0] fbank_1_temp;
    reg [31:0] fbank_2_temp;
    reg [31:0] fbank_3_temp;
    reg [31:0] fbank_4_temp;
    reg [31:0] fbank_5_temp;
    reg [31:0] fbank_6_temp;
    reg [31:0] fbank_7_temp;
    reg [31:0] fbank_8_temp;
    reg [31:0] fbank_9_temp;
    reg [31:0] fbank_10_temp;
    reg [31:0] fbank_11_temp;
    reg [31:0] fbank_12_temp;
    reg [31:0] fbank_13_temp;
    reg [31:0] fbank_14_temp;
    reg [31:0] fbank_15_temp;
    reg [31:0] fbank_16_temp;
    reg [31:0] fbank_17_temp;
    reg [31:0] fbank_18_temp;
    reg [31:0] fbank_19_temp;
    reg [31:0] fbank_20_temp;
    reg [31:0] fbank_21_temp;
    reg [31:0] fbank_22_temp;
    reg [31:0] fbank_23_temp;
    reg [31:0] fbank_24_temp;
    reg [31:0] fbank_25_temp;
    reg [31:0] fbank_26_temp;
    
    reg [4:0] cnt_feat = 0;
    
assign filter_banks_1[0] = 32'h00000000;
assign filter_banks_1[1] = 32'h3f000000;
assign filter_banks_1[2] = 32'h3f800000;
assign filter_banks_1[3] = 32'h3f000000;
assign filter_banks_1[4] = 32'h00000000;
assign filter_banks_1[5] = 32'h00000000;
assign filter_banks_1[6] = 32'h00000000;
assign filter_banks_1[7] = 32'h00000000;
assign filter_banks_1[8] = 32'h00000000;
assign filter_banks_1[9] = 32'h00000000;
assign filter_banks_1[10] = 32'h00000000;
assign filter_banks_1[11] = 32'h00000000;
assign filter_banks_1[12] = 32'h00000000;
assign filter_banks_1[13] = 32'h00000000;
assign filter_banks_1[14] = 32'h00000000;
assign filter_banks_1[15] = 32'h00000000;
assign filter_banks_1[16] = 32'h00000000;
assign filter_banks_1[17] = 32'h00000000;
assign filter_banks_1[18] = 32'h00000000;
assign filter_banks_1[19] = 32'h00000000;
assign filter_banks_1[20] = 32'h00000000;
assign filter_banks_1[21] = 32'h00000000;
assign filter_banks_1[22] = 32'h00000000;
assign filter_banks_1[23] = 32'h00000000;
assign filter_banks_1[24] = 32'h00000000;
assign filter_banks_1[25] = 32'h00000000;
assign filter_banks_1[26] = 32'h00000000;
assign filter_banks_1[27] = 32'h00000000;
assign filter_banks_1[28] = 32'h00000000;
assign filter_banks_1[29] = 32'h00000000;
assign filter_banks_1[30] = 32'h00000000;
assign filter_banks_1[31] = 32'h00000000;
assign filter_banks_1[32] = 32'h00000000;
assign filter_banks_1[33] = 32'h00000000;
assign filter_banks_1[34] = 32'h00000000;
assign filter_banks_1[35] = 32'h00000000;
assign filter_banks_1[36] = 32'h00000000;
assign filter_banks_1[37] = 32'h00000000;
assign filter_banks_1[38] = 32'h00000000;
assign filter_banks_1[39] = 32'h00000000;
assign filter_banks_1[40] = 32'h00000000;
assign filter_banks_1[41] = 32'h00000000;
assign filter_banks_1[42] = 32'h00000000;
assign filter_banks_1[43] = 32'h00000000;
assign filter_banks_1[44] = 32'h00000000;
assign filter_banks_1[45] = 32'h00000000;
assign filter_banks_1[46] = 32'h00000000;
assign filter_banks_1[47] = 32'h00000000;
assign filter_banks_1[48] = 32'h00000000;
assign filter_banks_1[49] = 32'h00000000;
assign filter_banks_1[50] = 32'h00000000;
assign filter_banks_1[51] = 32'h00000000;
assign filter_banks_1[52] = 32'h00000000;
assign filter_banks_1[53] = 32'h00000000;
assign filter_banks_1[54] = 32'h00000000;
assign filter_banks_1[55] = 32'h00000000;
assign filter_banks_1[56] = 32'h00000000;
assign filter_banks_1[57] = 32'h00000000;
assign filter_banks_1[58] = 32'h00000000;
assign filter_banks_1[59] = 32'h00000000;
assign filter_banks_1[60] = 32'h00000000;
assign filter_banks_1[61] = 32'h00000000;
assign filter_banks_1[62] = 32'h00000000;
assign filter_banks_1[63] = 32'h00000000;
assign filter_banks_1[64] = 32'h00000000;
assign filter_banks_1[65] = 32'h00000000;
assign filter_banks_1[66] = 32'h00000000;
assign filter_banks_1[67] = 32'h00000000;
assign filter_banks_1[68] = 32'h00000000;
assign filter_banks_1[69] = 32'h00000000;
assign filter_banks_1[70] = 32'h00000000;
assign filter_banks_1[71] = 32'h00000000;
assign filter_banks_1[72] = 32'h00000000;
assign filter_banks_1[73] = 32'h00000000;
assign filter_banks_1[74] = 32'h00000000;
assign filter_banks_1[75] = 32'h00000000;
assign filter_banks_1[76] = 32'h00000000;
assign filter_banks_1[77] = 32'h00000000;
assign filter_banks_1[78] = 32'h00000000;
assign filter_banks_1[79] = 32'h00000000;
assign filter_banks_1[80] = 32'h00000000;
assign filter_banks_1[81] = 32'h00000000;
assign filter_banks_1[82] = 32'h00000000;
assign filter_banks_1[83] = 32'h00000000;
assign filter_banks_1[84] = 32'h00000000;
assign filter_banks_1[85] = 32'h00000000;
assign filter_banks_1[86] = 32'h00000000;
assign filter_banks_1[87] = 32'h00000000;
assign filter_banks_1[88] = 32'h00000000;
assign filter_banks_1[89] = 32'h00000000;
assign filter_banks_1[90] = 32'h00000000;
assign filter_banks_1[91] = 32'h00000000;
assign filter_banks_1[92] = 32'h00000000;
assign filter_banks_1[93] = 32'h00000000;
assign filter_banks_1[94] = 32'h00000000;
assign filter_banks_1[95] = 32'h00000000;
assign filter_banks_1[96] = 32'h00000000;
assign filter_banks_1[97] = 32'h00000000;
assign filter_banks_1[98] = 32'h00000000;
assign filter_banks_1[99] = 32'h00000000;
assign filter_banks_1[100] = 32'h00000000;
assign filter_banks_1[101] = 32'h00000000;
assign filter_banks_1[102] = 32'h00000000;
assign filter_banks_1[103] = 32'h00000000;
assign filter_banks_1[104] = 32'h00000000;
assign filter_banks_1[105] = 32'h00000000;
assign filter_banks_1[106] = 32'h00000000;
assign filter_banks_1[107] = 32'h00000000;
assign filter_banks_1[108] = 32'h00000000;
assign filter_banks_1[109] = 32'h00000000;
assign filter_banks_1[110] = 32'h00000000;
assign filter_banks_1[111] = 32'h00000000;
assign filter_banks_1[112] = 32'h00000000;
assign filter_banks_1[113] = 32'h00000000;
assign filter_banks_1[114] = 32'h00000000;
assign filter_banks_1[115] = 32'h00000000;
assign filter_banks_1[116] = 32'h00000000;
assign filter_banks_1[117] = 32'h00000000;
assign filter_banks_1[118] = 32'h00000000;
assign filter_banks_1[119] = 32'h00000000;
assign filter_banks_1[120] = 32'h00000000;
assign filter_banks_1[121] = 32'h00000000;
assign filter_banks_1[122] = 32'h00000000;
assign filter_banks_1[123] = 32'h00000000;
assign filter_banks_1[124] = 32'h00000000;
assign filter_banks_1[125] = 32'h00000000;
assign filter_banks_1[126] = 32'h00000000;
assign filter_banks_1[127] = 32'h00000000;
assign filter_banks_1[128] = 32'h00000000;
assign filter_banks_1[129] = 32'h00000000;
assign filter_banks_1[130] = 32'h00000000;
assign filter_banks_1[131] = 32'h00000000;
assign filter_banks_1[132] = 32'h00000000;
assign filter_banks_1[133] = 32'h00000000;
assign filter_banks_1[134] = 32'h00000000;
assign filter_banks_1[135] = 32'h00000000;
assign filter_banks_1[136] = 32'h00000000;
assign filter_banks_1[137] = 32'h00000000;
assign filter_banks_1[138] = 32'h00000000;
assign filter_banks_1[139] = 32'h00000000;
assign filter_banks_1[140] = 32'h00000000;
assign filter_banks_1[141] = 32'h00000000;
assign filter_banks_1[142] = 32'h00000000;
assign filter_banks_1[143] = 32'h00000000;
assign filter_banks_1[144] = 32'h00000000;
assign filter_banks_1[145] = 32'h00000000;
assign filter_banks_1[146] = 32'h00000000;
assign filter_banks_1[147] = 32'h00000000;
assign filter_banks_1[148] = 32'h00000000;
assign filter_banks_1[149] = 32'h00000000;
assign filter_banks_1[150] = 32'h00000000;
assign filter_banks_1[151] = 32'h00000000;
assign filter_banks_1[152] = 32'h00000000;
assign filter_banks_1[153] = 32'h00000000;
assign filter_banks_1[154] = 32'h00000000;
assign filter_banks_1[155] = 32'h00000000;
assign filter_banks_1[156] = 32'h00000000;
assign filter_banks_1[157] = 32'h00000000;
assign filter_banks_1[158] = 32'h00000000;
assign filter_banks_1[159] = 32'h00000000;
assign filter_banks_1[160] = 32'h00000000;
assign filter_banks_1[161] = 32'h00000000;
assign filter_banks_1[162] = 32'h00000000;
assign filter_banks_1[163] = 32'h00000000;
assign filter_banks_1[164] = 32'h00000000;
assign filter_banks_1[165] = 32'h00000000;
assign filter_banks_1[166] = 32'h00000000;
assign filter_banks_1[167] = 32'h00000000;
assign filter_banks_1[168] = 32'h00000000;
assign filter_banks_1[169] = 32'h00000000;
assign filter_banks_1[170] = 32'h00000000;
assign filter_banks_1[171] = 32'h00000000;
assign filter_banks_1[172] = 32'h00000000;
assign filter_banks_1[173] = 32'h00000000;
assign filter_banks_1[174] = 32'h00000000;
assign filter_banks_1[175] = 32'h00000000;
assign filter_banks_1[176] = 32'h00000000;
assign filter_banks_1[177] = 32'h00000000;
assign filter_banks_1[178] = 32'h00000000;
assign filter_banks_1[179] = 32'h00000000;
assign filter_banks_1[180] = 32'h00000000;
assign filter_banks_1[181] = 32'h00000000;
assign filter_banks_1[182] = 32'h00000000;
assign filter_banks_1[183] = 32'h00000000;
assign filter_banks_1[184] = 32'h00000000;
assign filter_banks_1[185] = 32'h00000000;
assign filter_banks_1[186] = 32'h00000000;
assign filter_banks_1[187] = 32'h00000000;
assign filter_banks_1[188] = 32'h00000000;
assign filter_banks_1[189] = 32'h00000000;
assign filter_banks_1[190] = 32'h00000000;
assign filter_banks_1[191] = 32'h00000000;
assign filter_banks_1[192] = 32'h00000000;
assign filter_banks_1[193] = 32'h00000000;
assign filter_banks_1[194] = 32'h00000000;
assign filter_banks_1[195] = 32'h00000000;
assign filter_banks_1[196] = 32'h00000000;
assign filter_banks_1[197] = 32'h00000000;
assign filter_banks_1[198] = 32'h00000000;
assign filter_banks_1[199] = 32'h00000000;
assign filter_banks_1[200] = 32'h00000000;
assign filter_banks_1[201] = 32'h00000000;
assign filter_banks_1[202] = 32'h00000000;
assign filter_banks_1[203] = 32'h00000000;
assign filter_banks_1[204] = 32'h00000000;
assign filter_banks_1[205] = 32'h00000000;
assign filter_banks_1[206] = 32'h00000000;
assign filter_banks_1[207] = 32'h00000000;
assign filter_banks_1[208] = 32'h00000000;
assign filter_banks_1[209] = 32'h00000000;
assign filter_banks_1[210] = 32'h00000000;
assign filter_banks_1[211] = 32'h00000000;
assign filter_banks_1[212] = 32'h00000000;
assign filter_banks_1[213] = 32'h00000000;
assign filter_banks_1[214] = 32'h00000000;
assign filter_banks_1[215] = 32'h00000000;
assign filter_banks_1[216] = 32'h00000000;
assign filter_banks_1[217] = 32'h00000000;
assign filter_banks_1[218] = 32'h00000000;
assign filter_banks_1[219] = 32'h00000000;
assign filter_banks_1[220] = 32'h00000000;
assign filter_banks_1[221] = 32'h00000000;
assign filter_banks_1[222] = 32'h00000000;
assign filter_banks_1[223] = 32'h00000000;
assign filter_banks_1[224] = 32'h00000000;
assign filter_banks_1[225] = 32'h00000000;
assign filter_banks_1[226] = 32'h00000000;
assign filter_banks_1[227] = 32'h00000000;
assign filter_banks_1[228] = 32'h00000000;
assign filter_banks_1[229] = 32'h00000000;
assign filter_banks_1[230] = 32'h00000000;
assign filter_banks_1[231] = 32'h00000000;
assign filter_banks_1[232] = 32'h00000000;
assign filter_banks_1[233] = 32'h00000000;
assign filter_banks_1[234] = 32'h00000000;
assign filter_banks_1[235] = 32'h00000000;
assign filter_banks_1[236] = 32'h00000000;
assign filter_banks_1[237] = 32'h00000000;
assign filter_banks_1[238] = 32'h00000000;
assign filter_banks_1[239] = 32'h00000000;
assign filter_banks_1[240] = 32'h00000000;
assign filter_banks_1[241] = 32'h00000000;
assign filter_banks_1[242] = 32'h00000000;
assign filter_banks_1[243] = 32'h00000000;
assign filter_banks_1[244] = 32'h00000000;
assign filter_banks_1[245] = 32'h00000000;
assign filter_banks_1[246] = 32'h00000000;
assign filter_banks_1[247] = 32'h00000000;
assign filter_banks_1[248] = 32'h00000000;
assign filter_banks_1[249] = 32'h00000000;
assign filter_banks_1[250] = 32'h00000000;
assign filter_banks_1[251] = 32'h00000000;
assign filter_banks_1[252] = 32'h00000000;
assign filter_banks_1[253] = 32'h00000000;
assign filter_banks_1[254] = 32'h00000000;
assign filter_banks_1[255] = 32'h00000000;
assign filter_banks_1[256] = 32'h00000000;
assign filter_banks_2[0] = 32'h00000000;
assign filter_banks_2[1] = 32'h00000000;
assign filter_banks_2[2] = 32'h00000000;
assign filter_banks_2[3] = 32'h3f000000;
assign filter_banks_2[4] = 32'h3f800000;
assign filter_banks_2[5] = 32'h3f2aaaab;
assign filter_banks_2[6] = 32'h3eaaaaab;
assign filter_banks_2[7] = 32'h00000000;
assign filter_banks_2[8] = 32'h00000000;
assign filter_banks_2[9] = 32'h00000000;
assign filter_banks_2[10] = 32'h00000000;
assign filter_banks_2[11] = 32'h00000000;
assign filter_banks_2[12] = 32'h00000000;
assign filter_banks_2[13] = 32'h00000000;
assign filter_banks_2[14] = 32'h00000000;
assign filter_banks_2[15] = 32'h00000000;
assign filter_banks_2[16] = 32'h00000000;
assign filter_banks_2[17] = 32'h00000000;
assign filter_banks_2[18] = 32'h00000000;
assign filter_banks_2[19] = 32'h00000000;
assign filter_banks_2[20] = 32'h00000000;
assign filter_banks_2[21] = 32'h00000000;
assign filter_banks_2[22] = 32'h00000000;
assign filter_banks_2[23] = 32'h00000000;
assign filter_banks_2[24] = 32'h00000000;
assign filter_banks_2[25] = 32'h00000000;
assign filter_banks_2[26] = 32'h00000000;
assign filter_banks_2[27] = 32'h00000000;
assign filter_banks_2[28] = 32'h00000000;
assign filter_banks_2[29] = 32'h00000000;
assign filter_banks_2[30] = 32'h00000000;
assign filter_banks_2[31] = 32'h00000000;
assign filter_banks_2[32] = 32'h00000000;
assign filter_banks_2[33] = 32'h00000000;
assign filter_banks_2[34] = 32'h00000000;
assign filter_banks_2[35] = 32'h00000000;
assign filter_banks_2[36] = 32'h00000000;
assign filter_banks_2[37] = 32'h00000000;
assign filter_banks_2[38] = 32'h00000000;
assign filter_banks_2[39] = 32'h00000000;
assign filter_banks_2[40] = 32'h00000000;
assign filter_banks_2[41] = 32'h00000000;
assign filter_banks_2[42] = 32'h00000000;
assign filter_banks_2[43] = 32'h00000000;
assign filter_banks_2[44] = 32'h00000000;
assign filter_banks_2[45] = 32'h00000000;
assign filter_banks_2[46] = 32'h00000000;
assign filter_banks_2[47] = 32'h00000000;
assign filter_banks_2[48] = 32'h00000000;
assign filter_banks_2[49] = 32'h00000000;
assign filter_banks_2[50] = 32'h00000000;
assign filter_banks_2[51] = 32'h00000000;
assign filter_banks_2[52] = 32'h00000000;
assign filter_banks_2[53] = 32'h00000000;
assign filter_banks_2[54] = 32'h00000000;
assign filter_banks_2[55] = 32'h00000000;
assign filter_banks_2[56] = 32'h00000000;
assign filter_banks_2[57] = 32'h00000000;
assign filter_banks_2[58] = 32'h00000000;
assign filter_banks_2[59] = 32'h00000000;
assign filter_banks_2[60] = 32'h00000000;
assign filter_banks_2[61] = 32'h00000000;
assign filter_banks_2[62] = 32'h00000000;
assign filter_banks_2[63] = 32'h00000000;
assign filter_banks_2[64] = 32'h00000000;
assign filter_banks_2[65] = 32'h00000000;
assign filter_banks_2[66] = 32'h00000000;
assign filter_banks_2[67] = 32'h00000000;
assign filter_banks_2[68] = 32'h00000000;
assign filter_banks_2[69] = 32'h00000000;
assign filter_banks_2[70] = 32'h00000000;
assign filter_banks_2[71] = 32'h00000000;
assign filter_banks_2[72] = 32'h00000000;
assign filter_banks_2[73] = 32'h00000000;
assign filter_banks_2[74] = 32'h00000000;
assign filter_banks_2[75] = 32'h00000000;
assign filter_banks_2[76] = 32'h00000000;
assign filter_banks_2[77] = 32'h00000000;
assign filter_banks_2[78] = 32'h00000000;
assign filter_banks_2[79] = 32'h00000000;
assign filter_banks_2[80] = 32'h00000000;
assign filter_banks_2[81] = 32'h00000000;
assign filter_banks_2[82] = 32'h00000000;
assign filter_banks_2[83] = 32'h00000000;
assign filter_banks_2[84] = 32'h00000000;
assign filter_banks_2[85] = 32'h00000000;
assign filter_banks_2[86] = 32'h00000000;
assign filter_banks_2[87] = 32'h00000000;
assign filter_banks_2[88] = 32'h00000000;
assign filter_banks_2[89] = 32'h00000000;
assign filter_banks_2[90] = 32'h00000000;
assign filter_banks_2[91] = 32'h00000000;
assign filter_banks_2[92] = 32'h00000000;
assign filter_banks_2[93] = 32'h00000000;
assign filter_banks_2[94] = 32'h00000000;
assign filter_banks_2[95] = 32'h00000000;
assign filter_banks_2[96] = 32'h00000000;
assign filter_banks_2[97] = 32'h00000000;
assign filter_banks_2[98] = 32'h00000000;
assign filter_banks_2[99] = 32'h00000000;
assign filter_banks_2[100] = 32'h00000000;
assign filter_banks_2[101] = 32'h00000000;
assign filter_banks_2[102] = 32'h00000000;
assign filter_banks_2[103] = 32'h00000000;
assign filter_banks_2[104] = 32'h00000000;
assign filter_banks_2[105] = 32'h00000000;
assign filter_banks_2[106] = 32'h00000000;
assign filter_banks_2[107] = 32'h00000000;
assign filter_banks_2[108] = 32'h00000000;
assign filter_banks_2[109] = 32'h00000000;
assign filter_banks_2[110] = 32'h00000000;
assign filter_banks_2[111] = 32'h00000000;
assign filter_banks_2[112] = 32'h00000000;
assign filter_banks_2[113] = 32'h00000000;
assign filter_banks_2[114] = 32'h00000000;
assign filter_banks_2[115] = 32'h00000000;
assign filter_banks_2[116] = 32'h00000000;
assign filter_banks_2[117] = 32'h00000000;
assign filter_banks_2[118] = 32'h00000000;
assign filter_banks_2[119] = 32'h00000000;
assign filter_banks_2[120] = 32'h00000000;
assign filter_banks_2[121] = 32'h00000000;
assign filter_banks_2[122] = 32'h00000000;
assign filter_banks_2[123] = 32'h00000000;
assign filter_banks_2[124] = 32'h00000000;
assign filter_banks_2[125] = 32'h00000000;
assign filter_banks_2[126] = 32'h00000000;
assign filter_banks_2[127] = 32'h00000000;
assign filter_banks_2[128] = 32'h00000000;
assign filter_banks_2[129] = 32'h00000000;
assign filter_banks_2[130] = 32'h00000000;
assign filter_banks_2[131] = 32'h00000000;
assign filter_banks_2[132] = 32'h00000000;
assign filter_banks_2[133] = 32'h00000000;
assign filter_banks_2[134] = 32'h00000000;
assign filter_banks_2[135] = 32'h00000000;
assign filter_banks_2[136] = 32'h00000000;
assign filter_banks_2[137] = 32'h00000000;
assign filter_banks_2[138] = 32'h00000000;
assign filter_banks_2[139] = 32'h00000000;
assign filter_banks_2[140] = 32'h00000000;
assign filter_banks_2[141] = 32'h00000000;
assign filter_banks_2[142] = 32'h00000000;
assign filter_banks_2[143] = 32'h00000000;
assign filter_banks_2[144] = 32'h00000000;
assign filter_banks_2[145] = 32'h00000000;
assign filter_banks_2[146] = 32'h00000000;
assign filter_banks_2[147] = 32'h00000000;
assign filter_banks_2[148] = 32'h00000000;
assign filter_banks_2[149] = 32'h00000000;
assign filter_banks_2[150] = 32'h00000000;
assign filter_banks_2[151] = 32'h00000000;
assign filter_banks_2[152] = 32'h00000000;
assign filter_banks_2[153] = 32'h00000000;
assign filter_banks_2[154] = 32'h00000000;
assign filter_banks_2[155] = 32'h00000000;
assign filter_banks_2[156] = 32'h00000000;
assign filter_banks_2[157] = 32'h00000000;
assign filter_banks_2[158] = 32'h00000000;
assign filter_banks_2[159] = 32'h00000000;
assign filter_banks_2[160] = 32'h00000000;
assign filter_banks_2[161] = 32'h00000000;
assign filter_banks_2[162] = 32'h00000000;
assign filter_banks_2[163] = 32'h00000000;
assign filter_banks_2[164] = 32'h00000000;
assign filter_banks_2[165] = 32'h00000000;
assign filter_banks_2[166] = 32'h00000000;
assign filter_banks_2[167] = 32'h00000000;
assign filter_banks_2[168] = 32'h00000000;
assign filter_banks_2[169] = 32'h00000000;
assign filter_banks_2[170] = 32'h00000000;
assign filter_banks_2[171] = 32'h00000000;
assign filter_banks_2[172] = 32'h00000000;
assign filter_banks_2[173] = 32'h00000000;
assign filter_banks_2[174] = 32'h00000000;
assign filter_banks_2[175] = 32'h00000000;
assign filter_banks_2[176] = 32'h00000000;
assign filter_banks_2[177] = 32'h00000000;
assign filter_banks_2[178] = 32'h00000000;
assign filter_banks_2[179] = 32'h00000000;
assign filter_banks_2[180] = 32'h00000000;
assign filter_banks_2[181] = 32'h00000000;
assign filter_banks_2[182] = 32'h00000000;
assign filter_banks_2[183] = 32'h00000000;
assign filter_banks_2[184] = 32'h00000000;
assign filter_banks_2[185] = 32'h00000000;
assign filter_banks_2[186] = 32'h00000000;
assign filter_banks_2[187] = 32'h00000000;
assign filter_banks_2[188] = 32'h00000000;
assign filter_banks_2[189] = 32'h00000000;
assign filter_banks_2[190] = 32'h00000000;
assign filter_banks_2[191] = 32'h00000000;
assign filter_banks_2[192] = 32'h00000000;
assign filter_banks_2[193] = 32'h00000000;
assign filter_banks_2[194] = 32'h00000000;
assign filter_banks_2[195] = 32'h00000000;
assign filter_banks_2[196] = 32'h00000000;
assign filter_banks_2[197] = 32'h00000000;
assign filter_banks_2[198] = 32'h00000000;
assign filter_banks_2[199] = 32'h00000000;
assign filter_banks_2[200] = 32'h00000000;
assign filter_banks_2[201] = 32'h00000000;
assign filter_banks_2[202] = 32'h00000000;
assign filter_banks_2[203] = 32'h00000000;
assign filter_banks_2[204] = 32'h00000000;
assign filter_banks_2[205] = 32'h00000000;
assign filter_banks_2[206] = 32'h00000000;
assign filter_banks_2[207] = 32'h00000000;
assign filter_banks_2[208] = 32'h00000000;
assign filter_banks_2[209] = 32'h00000000;
assign filter_banks_2[210] = 32'h00000000;
assign filter_banks_2[211] = 32'h00000000;
assign filter_banks_2[212] = 32'h00000000;
assign filter_banks_2[213] = 32'h00000000;
assign filter_banks_2[214] = 32'h00000000;
assign filter_banks_2[215] = 32'h00000000;
assign filter_banks_2[216] = 32'h00000000;
assign filter_banks_2[217] = 32'h00000000;
assign filter_banks_2[218] = 32'h00000000;
assign filter_banks_2[219] = 32'h00000000;
assign filter_banks_2[220] = 32'h00000000;
assign filter_banks_2[221] = 32'h00000000;
assign filter_banks_2[222] = 32'h00000000;
assign filter_banks_2[223] = 32'h00000000;
assign filter_banks_2[224] = 32'h00000000;
assign filter_banks_2[225] = 32'h00000000;
assign filter_banks_2[226] = 32'h00000000;
assign filter_banks_2[227] = 32'h00000000;
assign filter_banks_2[228] = 32'h00000000;
assign filter_banks_2[229] = 32'h00000000;
assign filter_banks_2[230] = 32'h00000000;
assign filter_banks_2[231] = 32'h00000000;
assign filter_banks_2[232] = 32'h00000000;
assign filter_banks_2[233] = 32'h00000000;
assign filter_banks_2[234] = 32'h00000000;
assign filter_banks_2[235] = 32'h00000000;
assign filter_banks_2[236] = 32'h00000000;
assign filter_banks_2[237] = 32'h00000000;
assign filter_banks_2[238] = 32'h00000000;
assign filter_banks_2[239] = 32'h00000000;
assign filter_banks_2[240] = 32'h00000000;
assign filter_banks_2[241] = 32'h00000000;
assign filter_banks_2[242] = 32'h00000000;
assign filter_banks_2[243] = 32'h00000000;
assign filter_banks_2[244] = 32'h00000000;
assign filter_banks_2[245] = 32'h00000000;
assign filter_banks_2[246] = 32'h00000000;
assign filter_banks_2[247] = 32'h00000000;
assign filter_banks_2[248] = 32'h00000000;
assign filter_banks_2[249] = 32'h00000000;
assign filter_banks_2[250] = 32'h00000000;
assign filter_banks_2[251] = 32'h00000000;
assign filter_banks_2[252] = 32'h00000000;
assign filter_banks_2[253] = 32'h00000000;
assign filter_banks_2[254] = 32'h00000000;
assign filter_banks_2[255] = 32'h00000000;
assign filter_banks_2[256] = 32'h00000000;
assign filter_banks_3[0] = 32'h00000000;
assign filter_banks_3[1] = 32'h00000000;
assign filter_banks_3[2] = 32'h00000000;
assign filter_banks_3[3] = 32'h00000000;
assign filter_banks_3[4] = 32'h00000000;
assign filter_banks_3[5] = 32'h3eaaaaab;
assign filter_banks_3[6] = 32'h3f2aaaab;
assign filter_banks_3[7] = 32'h3f800000;
assign filter_banks_3[8] = 32'h3f2aaaab;
assign filter_banks_3[9] = 32'h3eaaaaab;
assign filter_banks_3[10] = 32'h00000000;
assign filter_banks_3[11] = 32'h00000000;
assign filter_banks_3[12] = 32'h00000000;
assign filter_banks_3[13] = 32'h00000000;
assign filter_banks_3[14] = 32'h00000000;
assign filter_banks_3[15] = 32'h00000000;
assign filter_banks_3[16] = 32'h00000000;
assign filter_banks_3[17] = 32'h00000000;
assign filter_banks_3[18] = 32'h00000000;
assign filter_banks_3[19] = 32'h00000000;
assign filter_banks_3[20] = 32'h00000000;
assign filter_banks_3[21] = 32'h00000000;
assign filter_banks_3[22] = 32'h00000000;
assign filter_banks_3[23] = 32'h00000000;
assign filter_banks_3[24] = 32'h00000000;
assign filter_banks_3[25] = 32'h00000000;
assign filter_banks_3[26] = 32'h00000000;
assign filter_banks_3[27] = 32'h00000000;
assign filter_banks_3[28] = 32'h00000000;
assign filter_banks_3[29] = 32'h00000000;
assign filter_banks_3[30] = 32'h00000000;
assign filter_banks_3[31] = 32'h00000000;
assign filter_banks_3[32] = 32'h00000000;
assign filter_banks_3[33] = 32'h00000000;
assign filter_banks_3[34] = 32'h00000000;
assign filter_banks_3[35] = 32'h00000000;
assign filter_banks_3[36] = 32'h00000000;
assign filter_banks_3[37] = 32'h00000000;
assign filter_banks_3[38] = 32'h00000000;
assign filter_banks_3[39] = 32'h00000000;
assign filter_banks_3[40] = 32'h00000000;
assign filter_banks_3[41] = 32'h00000000;
assign filter_banks_3[42] = 32'h00000000;
assign filter_banks_3[43] = 32'h00000000;
assign filter_banks_3[44] = 32'h00000000;
assign filter_banks_3[45] = 32'h00000000;
assign filter_banks_3[46] = 32'h00000000;
assign filter_banks_3[47] = 32'h00000000;
assign filter_banks_3[48] = 32'h00000000;
assign filter_banks_3[49] = 32'h00000000;
assign filter_banks_3[50] = 32'h00000000;
assign filter_banks_3[51] = 32'h00000000;
assign filter_banks_3[52] = 32'h00000000;
assign filter_banks_3[53] = 32'h00000000;
assign filter_banks_3[54] = 32'h00000000;
assign filter_banks_3[55] = 32'h00000000;
assign filter_banks_3[56] = 32'h00000000;
assign filter_banks_3[57] = 32'h00000000;
assign filter_banks_3[58] = 32'h00000000;
assign filter_banks_3[59] = 32'h00000000;
assign filter_banks_3[60] = 32'h00000000;
assign filter_banks_3[61] = 32'h00000000;
assign filter_banks_3[62] = 32'h00000000;
assign filter_banks_3[63] = 32'h00000000;
assign filter_banks_3[64] = 32'h00000000;
assign filter_banks_3[65] = 32'h00000000;
assign filter_banks_3[66] = 32'h00000000;
assign filter_banks_3[67] = 32'h00000000;
assign filter_banks_3[68] = 32'h00000000;
assign filter_banks_3[69] = 32'h00000000;
assign filter_banks_3[70] = 32'h00000000;
assign filter_banks_3[71] = 32'h00000000;
assign filter_banks_3[72] = 32'h00000000;
assign filter_banks_3[73] = 32'h00000000;
assign filter_banks_3[74] = 32'h00000000;
assign filter_banks_3[75] = 32'h00000000;
assign filter_banks_3[76] = 32'h00000000;
assign filter_banks_3[77] = 32'h00000000;
assign filter_banks_3[78] = 32'h00000000;
assign filter_banks_3[79] = 32'h00000000;
assign filter_banks_3[80] = 32'h00000000;
assign filter_banks_3[81] = 32'h00000000;
assign filter_banks_3[82] = 32'h00000000;
assign filter_banks_3[83] = 32'h00000000;
assign filter_banks_3[84] = 32'h00000000;
assign filter_banks_3[85] = 32'h00000000;
assign filter_banks_3[86] = 32'h00000000;
assign filter_banks_3[87] = 32'h00000000;
assign filter_banks_3[88] = 32'h00000000;
assign filter_banks_3[89] = 32'h00000000;
assign filter_banks_3[90] = 32'h00000000;
assign filter_banks_3[91] = 32'h00000000;
assign filter_banks_3[92] = 32'h00000000;
assign filter_banks_3[93] = 32'h00000000;
assign filter_banks_3[94] = 32'h00000000;
assign filter_banks_3[95] = 32'h00000000;
assign filter_banks_3[96] = 32'h00000000;
assign filter_banks_3[97] = 32'h00000000;
assign filter_banks_3[98] = 32'h00000000;
assign filter_banks_3[99] = 32'h00000000;
assign filter_banks_3[100] = 32'h00000000;
assign filter_banks_3[101] = 32'h00000000;
assign filter_banks_3[102] = 32'h00000000;
assign filter_banks_3[103] = 32'h00000000;
assign filter_banks_3[104] = 32'h00000000;
assign filter_banks_3[105] = 32'h00000000;
assign filter_banks_3[106] = 32'h00000000;
assign filter_banks_3[107] = 32'h00000000;
assign filter_banks_3[108] = 32'h00000000;
assign filter_banks_3[109] = 32'h00000000;
assign filter_banks_3[110] = 32'h00000000;
assign filter_banks_3[111] = 32'h00000000;
assign filter_banks_3[112] = 32'h00000000;
assign filter_banks_3[113] = 32'h00000000;
assign filter_banks_3[114] = 32'h00000000;
assign filter_banks_3[115] = 32'h00000000;
assign filter_banks_3[116] = 32'h00000000;
assign filter_banks_3[117] = 32'h00000000;
assign filter_banks_3[118] = 32'h00000000;
assign filter_banks_3[119] = 32'h00000000;
assign filter_banks_3[120] = 32'h00000000;
assign filter_banks_3[121] = 32'h00000000;
assign filter_banks_3[122] = 32'h00000000;
assign filter_banks_3[123] = 32'h00000000;
assign filter_banks_3[124] = 32'h00000000;
assign filter_banks_3[125] = 32'h00000000;
assign filter_banks_3[126] = 32'h00000000;
assign filter_banks_3[127] = 32'h00000000;
assign filter_banks_3[128] = 32'h00000000;
assign filter_banks_3[129] = 32'h00000000;
assign filter_banks_3[130] = 32'h00000000;
assign filter_banks_3[131] = 32'h00000000;
assign filter_banks_3[132] = 32'h00000000;
assign filter_banks_3[133] = 32'h00000000;
assign filter_banks_3[134] = 32'h00000000;
assign filter_banks_3[135] = 32'h00000000;
assign filter_banks_3[136] = 32'h00000000;
assign filter_banks_3[137] = 32'h00000000;
assign filter_banks_3[138] = 32'h00000000;
assign filter_banks_3[139] = 32'h00000000;
assign filter_banks_3[140] = 32'h00000000;
assign filter_banks_3[141] = 32'h00000000;
assign filter_banks_3[142] = 32'h00000000;
assign filter_banks_3[143] = 32'h00000000;
assign filter_banks_3[144] = 32'h00000000;
assign filter_banks_3[145] = 32'h00000000;
assign filter_banks_3[146] = 32'h00000000;
assign filter_banks_3[147] = 32'h00000000;
assign filter_banks_3[148] = 32'h00000000;
assign filter_banks_3[149] = 32'h00000000;
assign filter_banks_3[150] = 32'h00000000;
assign filter_banks_3[151] = 32'h00000000;
assign filter_banks_3[152] = 32'h00000000;
assign filter_banks_3[153] = 32'h00000000;
assign filter_banks_3[154] = 32'h00000000;
assign filter_banks_3[155] = 32'h00000000;
assign filter_banks_3[156] = 32'h00000000;
assign filter_banks_3[157] = 32'h00000000;
assign filter_banks_3[158] = 32'h00000000;
assign filter_banks_3[159] = 32'h00000000;
assign filter_banks_3[160] = 32'h00000000;
assign filter_banks_3[161] = 32'h00000000;
assign filter_banks_3[162] = 32'h00000000;
assign filter_banks_3[163] = 32'h00000000;
assign filter_banks_3[164] = 32'h00000000;
assign filter_banks_3[165] = 32'h00000000;
assign filter_banks_3[166] = 32'h00000000;
assign filter_banks_3[167] = 32'h00000000;
assign filter_banks_3[168] = 32'h00000000;
assign filter_banks_3[169] = 32'h00000000;
assign filter_banks_3[170] = 32'h00000000;
assign filter_banks_3[171] = 32'h00000000;
assign filter_banks_3[172] = 32'h00000000;
assign filter_banks_3[173] = 32'h00000000;
assign filter_banks_3[174] = 32'h00000000;
assign filter_banks_3[175] = 32'h00000000;
assign filter_banks_3[176] = 32'h00000000;
assign filter_banks_3[177] = 32'h00000000;
assign filter_banks_3[178] = 32'h00000000;
assign filter_banks_3[179] = 32'h00000000;
assign filter_banks_3[180] = 32'h00000000;
assign filter_banks_3[181] = 32'h00000000;
assign filter_banks_3[182] = 32'h00000000;
assign filter_banks_3[183] = 32'h00000000;
assign filter_banks_3[184] = 32'h00000000;
assign filter_banks_3[185] = 32'h00000000;
assign filter_banks_3[186] = 32'h00000000;
assign filter_banks_3[187] = 32'h00000000;
assign filter_banks_3[188] = 32'h00000000;
assign filter_banks_3[189] = 32'h00000000;
assign filter_banks_3[190] = 32'h00000000;
assign filter_banks_3[191] = 32'h00000000;
assign filter_banks_3[192] = 32'h00000000;
assign filter_banks_3[193] = 32'h00000000;
assign filter_banks_3[194] = 32'h00000000;
assign filter_banks_3[195] = 32'h00000000;
assign filter_banks_3[196] = 32'h00000000;
assign filter_banks_3[197] = 32'h00000000;
assign filter_banks_3[198] = 32'h00000000;
assign filter_banks_3[199] = 32'h00000000;
assign filter_banks_3[200] = 32'h00000000;
assign filter_banks_3[201] = 32'h00000000;
assign filter_banks_3[202] = 32'h00000000;
assign filter_banks_3[203] = 32'h00000000;
assign filter_banks_3[204] = 32'h00000000;
assign filter_banks_3[205] = 32'h00000000;
assign filter_banks_3[206] = 32'h00000000;
assign filter_banks_3[207] = 32'h00000000;
assign filter_banks_3[208] = 32'h00000000;
assign filter_banks_3[209] = 32'h00000000;
assign filter_banks_3[210] = 32'h00000000;
assign filter_banks_3[211] = 32'h00000000;
assign filter_banks_3[212] = 32'h00000000;
assign filter_banks_3[213] = 32'h00000000;
assign filter_banks_3[214] = 32'h00000000;
assign filter_banks_3[215] = 32'h00000000;
assign filter_banks_3[216] = 32'h00000000;
assign filter_banks_3[217] = 32'h00000000;
assign filter_banks_3[218] = 32'h00000000;
assign filter_banks_3[219] = 32'h00000000;
assign filter_banks_3[220] = 32'h00000000;
assign filter_banks_3[221] = 32'h00000000;
assign filter_banks_3[222] = 32'h00000000;
assign filter_banks_3[223] = 32'h00000000;
assign filter_banks_3[224] = 32'h00000000;
assign filter_banks_3[225] = 32'h00000000;
assign filter_banks_3[226] = 32'h00000000;
assign filter_banks_3[227] = 32'h00000000;
assign filter_banks_3[228] = 32'h00000000;
assign filter_banks_3[229] = 32'h00000000;
assign filter_banks_3[230] = 32'h00000000;
assign filter_banks_3[231] = 32'h00000000;
assign filter_banks_3[232] = 32'h00000000;
assign filter_banks_3[233] = 32'h00000000;
assign filter_banks_3[234] = 32'h00000000;
assign filter_banks_3[235] = 32'h00000000;
assign filter_banks_3[236] = 32'h00000000;
assign filter_banks_3[237] = 32'h00000000;
assign filter_banks_3[238] = 32'h00000000;
assign filter_banks_3[239] = 32'h00000000;
assign filter_banks_3[240] = 32'h00000000;
assign filter_banks_3[241] = 32'h00000000;
assign filter_banks_3[242] = 32'h00000000;
assign filter_banks_3[243] = 32'h00000000;
assign filter_banks_3[244] = 32'h00000000;
assign filter_banks_3[245] = 32'h00000000;
assign filter_banks_3[246] = 32'h00000000;
assign filter_banks_3[247] = 32'h00000000;
assign filter_banks_3[248] = 32'h00000000;
assign filter_banks_3[249] = 32'h00000000;
assign filter_banks_3[250] = 32'h00000000;
assign filter_banks_3[251] = 32'h00000000;
assign filter_banks_3[252] = 32'h00000000;
assign filter_banks_3[253] = 32'h00000000;
assign filter_banks_3[254] = 32'h00000000;
assign filter_banks_3[255] = 32'h00000000;
assign filter_banks_3[256] = 32'h00000000;
assign filter_banks_4[0] = 32'h00000000;
assign filter_banks_4[1] = 32'h00000000;
assign filter_banks_4[2] = 32'h00000000;
assign filter_banks_4[3] = 32'h00000000;
assign filter_banks_4[4] = 32'h00000000;
assign filter_banks_4[5] = 32'h00000000;
assign filter_banks_4[6] = 32'h00000000;
assign filter_banks_4[7] = 32'h00000000;
assign filter_banks_4[8] = 32'h3eaaaaab;
assign filter_banks_4[9] = 32'h3f2aaaab;
assign filter_banks_4[10] = 32'h3f800000;
assign filter_banks_4[11] = 32'h3f2aaaab;
assign filter_banks_4[12] = 32'h3eaaaaab;
assign filter_banks_4[13] = 32'h00000000;
assign filter_banks_4[14] = 32'h00000000;
assign filter_banks_4[15] = 32'h00000000;
assign filter_banks_4[16] = 32'h00000000;
assign filter_banks_4[17] = 32'h00000000;
assign filter_banks_4[18] = 32'h00000000;
assign filter_banks_4[19] = 32'h00000000;
assign filter_banks_4[20] = 32'h00000000;
assign filter_banks_4[21] = 32'h00000000;
assign filter_banks_4[22] = 32'h00000000;
assign filter_banks_4[23] = 32'h00000000;
assign filter_banks_4[24] = 32'h00000000;
assign filter_banks_4[25] = 32'h00000000;
assign filter_banks_4[26] = 32'h00000000;
assign filter_banks_4[27] = 32'h00000000;
assign filter_banks_4[28] = 32'h00000000;
assign filter_banks_4[29] = 32'h00000000;
assign filter_banks_4[30] = 32'h00000000;
assign filter_banks_4[31] = 32'h00000000;
assign filter_banks_4[32] = 32'h00000000;
assign filter_banks_4[33] = 32'h00000000;
assign filter_banks_4[34] = 32'h00000000;
assign filter_banks_4[35] = 32'h00000000;
assign filter_banks_4[36] = 32'h00000000;
assign filter_banks_4[37] = 32'h00000000;
assign filter_banks_4[38] = 32'h00000000;
assign filter_banks_4[39] = 32'h00000000;
assign filter_banks_4[40] = 32'h00000000;
assign filter_banks_4[41] = 32'h00000000;
assign filter_banks_4[42] = 32'h00000000;
assign filter_banks_4[43] = 32'h00000000;
assign filter_banks_4[44] = 32'h00000000;
assign filter_banks_4[45] = 32'h00000000;
assign filter_banks_4[46] = 32'h00000000;
assign filter_banks_4[47] = 32'h00000000;
assign filter_banks_4[48] = 32'h00000000;
assign filter_banks_4[49] = 32'h00000000;
assign filter_banks_4[50] = 32'h00000000;
assign filter_banks_4[51] = 32'h00000000;
assign filter_banks_4[52] = 32'h00000000;
assign filter_banks_4[53] = 32'h00000000;
assign filter_banks_4[54] = 32'h00000000;
assign filter_banks_4[55] = 32'h00000000;
assign filter_banks_4[56] = 32'h00000000;
assign filter_banks_4[57] = 32'h00000000;
assign filter_banks_4[58] = 32'h00000000;
assign filter_banks_4[59] = 32'h00000000;
assign filter_banks_4[60] = 32'h00000000;
assign filter_banks_4[61] = 32'h00000000;
assign filter_banks_4[62] = 32'h00000000;
assign filter_banks_4[63] = 32'h00000000;
assign filter_banks_4[64] = 32'h00000000;
assign filter_banks_4[65] = 32'h00000000;
assign filter_banks_4[66] = 32'h00000000;
assign filter_banks_4[67] = 32'h00000000;
assign filter_banks_4[68] = 32'h00000000;
assign filter_banks_4[69] = 32'h00000000;
assign filter_banks_4[70] = 32'h00000000;
assign filter_banks_4[71] = 32'h00000000;
assign filter_banks_4[72] = 32'h00000000;
assign filter_banks_4[73] = 32'h00000000;
assign filter_banks_4[74] = 32'h00000000;
assign filter_banks_4[75] = 32'h00000000;
assign filter_banks_4[76] = 32'h00000000;
assign filter_banks_4[77] = 32'h00000000;
assign filter_banks_4[78] = 32'h00000000;
assign filter_banks_4[79] = 32'h00000000;
assign filter_banks_4[80] = 32'h00000000;
assign filter_banks_4[81] = 32'h00000000;
assign filter_banks_4[82] = 32'h00000000;
assign filter_banks_4[83] = 32'h00000000;
assign filter_banks_4[84] = 32'h00000000;
assign filter_banks_4[85] = 32'h00000000;
assign filter_banks_4[86] = 32'h00000000;
assign filter_banks_4[87] = 32'h00000000;
assign filter_banks_4[88] = 32'h00000000;
assign filter_banks_4[89] = 32'h00000000;
assign filter_banks_4[90] = 32'h00000000;
assign filter_banks_4[91] = 32'h00000000;
assign filter_banks_4[92] = 32'h00000000;
assign filter_banks_4[93] = 32'h00000000;
assign filter_banks_4[94] = 32'h00000000;
assign filter_banks_4[95] = 32'h00000000;
assign filter_banks_4[96] = 32'h00000000;
assign filter_banks_4[97] = 32'h00000000;
assign filter_banks_4[98] = 32'h00000000;
assign filter_banks_4[99] = 32'h00000000;
assign filter_banks_4[100] = 32'h00000000;
assign filter_banks_4[101] = 32'h00000000;
assign filter_banks_4[102] = 32'h00000000;
assign filter_banks_4[103] = 32'h00000000;
assign filter_banks_4[104] = 32'h00000000;
assign filter_banks_4[105] = 32'h00000000;
assign filter_banks_4[106] = 32'h00000000;
assign filter_banks_4[107] = 32'h00000000;
assign filter_banks_4[108] = 32'h00000000;
assign filter_banks_4[109] = 32'h00000000;
assign filter_banks_4[110] = 32'h00000000;
assign filter_banks_4[111] = 32'h00000000;
assign filter_banks_4[112] = 32'h00000000;
assign filter_banks_4[113] = 32'h00000000;
assign filter_banks_4[114] = 32'h00000000;
assign filter_banks_4[115] = 32'h00000000;
assign filter_banks_4[116] = 32'h00000000;
assign filter_banks_4[117] = 32'h00000000;
assign filter_banks_4[118] = 32'h00000000;
assign filter_banks_4[119] = 32'h00000000;
assign filter_banks_4[120] = 32'h00000000;
assign filter_banks_4[121] = 32'h00000000;
assign filter_banks_4[122] = 32'h00000000;
assign filter_banks_4[123] = 32'h00000000;
assign filter_banks_4[124] = 32'h00000000;
assign filter_banks_4[125] = 32'h00000000;
assign filter_banks_4[126] = 32'h00000000;
assign filter_banks_4[127] = 32'h00000000;
assign filter_banks_4[128] = 32'h00000000;
assign filter_banks_4[129] = 32'h00000000;
assign filter_banks_4[130] = 32'h00000000;
assign filter_banks_4[131] = 32'h00000000;
assign filter_banks_4[132] = 32'h00000000;
assign filter_banks_4[133] = 32'h00000000;
assign filter_banks_4[134] = 32'h00000000;
assign filter_banks_4[135] = 32'h00000000;
assign filter_banks_4[136] = 32'h00000000;
assign filter_banks_4[137] = 32'h00000000;
assign filter_banks_4[138] = 32'h00000000;
assign filter_banks_4[139] = 32'h00000000;
assign filter_banks_4[140] = 32'h00000000;
assign filter_banks_4[141] = 32'h00000000;
assign filter_banks_4[142] = 32'h00000000;
assign filter_banks_4[143] = 32'h00000000;
assign filter_banks_4[144] = 32'h00000000;
assign filter_banks_4[145] = 32'h00000000;
assign filter_banks_4[146] = 32'h00000000;
assign filter_banks_4[147] = 32'h00000000;
assign filter_banks_4[148] = 32'h00000000;
assign filter_banks_4[149] = 32'h00000000;
assign filter_banks_4[150] = 32'h00000000;
assign filter_banks_4[151] = 32'h00000000;
assign filter_banks_4[152] = 32'h00000000;
assign filter_banks_4[153] = 32'h00000000;
assign filter_banks_4[154] = 32'h00000000;
assign filter_banks_4[155] = 32'h00000000;
assign filter_banks_4[156] = 32'h00000000;
assign filter_banks_4[157] = 32'h00000000;
assign filter_banks_4[158] = 32'h00000000;
assign filter_banks_4[159] = 32'h00000000;
assign filter_banks_4[160] = 32'h00000000;
assign filter_banks_4[161] = 32'h00000000;
assign filter_banks_4[162] = 32'h00000000;
assign filter_banks_4[163] = 32'h00000000;
assign filter_banks_4[164] = 32'h00000000;
assign filter_banks_4[165] = 32'h00000000;
assign filter_banks_4[166] = 32'h00000000;
assign filter_banks_4[167] = 32'h00000000;
assign filter_banks_4[168] = 32'h00000000;
assign filter_banks_4[169] = 32'h00000000;
assign filter_banks_4[170] = 32'h00000000;
assign filter_banks_4[171] = 32'h00000000;
assign filter_banks_4[172] = 32'h00000000;
assign filter_banks_4[173] = 32'h00000000;
assign filter_banks_4[174] = 32'h00000000;
assign filter_banks_4[175] = 32'h00000000;
assign filter_banks_4[176] = 32'h00000000;
assign filter_banks_4[177] = 32'h00000000;
assign filter_banks_4[178] = 32'h00000000;
assign filter_banks_4[179] = 32'h00000000;
assign filter_banks_4[180] = 32'h00000000;
assign filter_banks_4[181] = 32'h00000000;
assign filter_banks_4[182] = 32'h00000000;
assign filter_banks_4[183] = 32'h00000000;
assign filter_banks_4[184] = 32'h00000000;
assign filter_banks_4[185] = 32'h00000000;
assign filter_banks_4[186] = 32'h00000000;
assign filter_banks_4[187] = 32'h00000000;
assign filter_banks_4[188] = 32'h00000000;
assign filter_banks_4[189] = 32'h00000000;
assign filter_banks_4[190] = 32'h00000000;
assign filter_banks_4[191] = 32'h00000000;
assign filter_banks_4[192] = 32'h00000000;
assign filter_banks_4[193] = 32'h00000000;
assign filter_banks_4[194] = 32'h00000000;
assign filter_banks_4[195] = 32'h00000000;
assign filter_banks_4[196] = 32'h00000000;
assign filter_banks_4[197] = 32'h00000000;
assign filter_banks_4[198] = 32'h00000000;
assign filter_banks_4[199] = 32'h00000000;
assign filter_banks_4[200] = 32'h00000000;
assign filter_banks_4[201] = 32'h00000000;
assign filter_banks_4[202] = 32'h00000000;
assign filter_banks_4[203] = 32'h00000000;
assign filter_banks_4[204] = 32'h00000000;
assign filter_banks_4[205] = 32'h00000000;
assign filter_banks_4[206] = 32'h00000000;
assign filter_banks_4[207] = 32'h00000000;
assign filter_banks_4[208] = 32'h00000000;
assign filter_banks_4[209] = 32'h00000000;
assign filter_banks_4[210] = 32'h00000000;
assign filter_banks_4[211] = 32'h00000000;
assign filter_banks_4[212] = 32'h00000000;
assign filter_banks_4[213] = 32'h00000000;
assign filter_banks_4[214] = 32'h00000000;
assign filter_banks_4[215] = 32'h00000000;
assign filter_banks_4[216] = 32'h00000000;
assign filter_banks_4[217] = 32'h00000000;
assign filter_banks_4[218] = 32'h00000000;
assign filter_banks_4[219] = 32'h00000000;
assign filter_banks_4[220] = 32'h00000000;
assign filter_banks_4[221] = 32'h00000000;
assign filter_banks_4[222] = 32'h00000000;
assign filter_banks_4[223] = 32'h00000000;
assign filter_banks_4[224] = 32'h00000000;
assign filter_banks_4[225] = 32'h00000000;
assign filter_banks_4[226] = 32'h00000000;
assign filter_banks_4[227] = 32'h00000000;
assign filter_banks_4[228] = 32'h00000000;
assign filter_banks_4[229] = 32'h00000000;
assign filter_banks_4[230] = 32'h00000000;
assign filter_banks_4[231] = 32'h00000000;
assign filter_banks_4[232] = 32'h00000000;
assign filter_banks_4[233] = 32'h00000000;
assign filter_banks_4[234] = 32'h00000000;
assign filter_banks_4[235] = 32'h00000000;
assign filter_banks_4[236] = 32'h00000000;
assign filter_banks_4[237] = 32'h00000000;
assign filter_banks_4[238] = 32'h00000000;
assign filter_banks_4[239] = 32'h00000000;
assign filter_banks_4[240] = 32'h00000000;
assign filter_banks_4[241] = 32'h00000000;
assign filter_banks_4[242] = 32'h00000000;
assign filter_banks_4[243] = 32'h00000000;
assign filter_banks_4[244] = 32'h00000000;
assign filter_banks_4[245] = 32'h00000000;
assign filter_banks_4[246] = 32'h00000000;
assign filter_banks_4[247] = 32'h00000000;
assign filter_banks_4[248] = 32'h00000000;
assign filter_banks_4[249] = 32'h00000000;
assign filter_banks_4[250] = 32'h00000000;
assign filter_banks_4[251] = 32'h00000000;
assign filter_banks_4[252] = 32'h00000000;
assign filter_banks_4[253] = 32'h00000000;
assign filter_banks_4[254] = 32'h00000000;
assign filter_banks_4[255] = 32'h00000000;
assign filter_banks_4[256] = 32'h00000000;
assign filter_banks_5[0] = 32'h00000000;
assign filter_banks_5[1] = 32'h00000000;
assign filter_banks_5[2] = 32'h00000000;
assign filter_banks_5[3] = 32'h00000000;
assign filter_banks_5[4] = 32'h00000000;
assign filter_banks_5[5] = 32'h00000000;
assign filter_banks_5[6] = 32'h00000000;
assign filter_banks_5[7] = 32'h00000000;
assign filter_banks_5[8] = 32'h00000000;
assign filter_banks_5[9] = 32'h00000000;
assign filter_banks_5[10] = 32'h00000000;
assign filter_banks_5[11] = 32'h3eaaaaab;
assign filter_banks_5[12] = 32'h3f2aaaab;
assign filter_banks_5[13] = 32'h3f800000;
assign filter_banks_5[14] = 32'h3f2aaaab;
assign filter_banks_5[15] = 32'h3eaaaaab;
assign filter_banks_5[16] = 32'h00000000;
assign filter_banks_5[17] = 32'h00000000;
assign filter_banks_5[18] = 32'h00000000;
assign filter_banks_5[19] = 32'h00000000;
assign filter_banks_5[20] = 32'h00000000;
assign filter_banks_5[21] = 32'h00000000;
assign filter_banks_5[22] = 32'h00000000;
assign filter_banks_5[23] = 32'h00000000;
assign filter_banks_5[24] = 32'h00000000;
assign filter_banks_5[25] = 32'h00000000;
assign filter_banks_5[26] = 32'h00000000;
assign filter_banks_5[27] = 32'h00000000;
assign filter_banks_5[28] = 32'h00000000;
assign filter_banks_5[29] = 32'h00000000;
assign filter_banks_5[30] = 32'h00000000;
assign filter_banks_5[31] = 32'h00000000;
assign filter_banks_5[32] = 32'h00000000;
assign filter_banks_5[33] = 32'h00000000;
assign filter_banks_5[34] = 32'h00000000;
assign filter_banks_5[35] = 32'h00000000;
assign filter_banks_5[36] = 32'h00000000;
assign filter_banks_5[37] = 32'h00000000;
assign filter_banks_5[38] = 32'h00000000;
assign filter_banks_5[39] = 32'h00000000;
assign filter_banks_5[40] = 32'h00000000;
assign filter_banks_5[41] = 32'h00000000;
assign filter_banks_5[42] = 32'h00000000;
assign filter_banks_5[43] = 32'h00000000;
assign filter_banks_5[44] = 32'h00000000;
assign filter_banks_5[45] = 32'h00000000;
assign filter_banks_5[46] = 32'h00000000;
assign filter_banks_5[47] = 32'h00000000;
assign filter_banks_5[48] = 32'h00000000;
assign filter_banks_5[49] = 32'h00000000;
assign filter_banks_5[50] = 32'h00000000;
assign filter_banks_5[51] = 32'h00000000;
assign filter_banks_5[52] = 32'h00000000;
assign filter_banks_5[53] = 32'h00000000;
assign filter_banks_5[54] = 32'h00000000;
assign filter_banks_5[55] = 32'h00000000;
assign filter_banks_5[56] = 32'h00000000;
assign filter_banks_5[57] = 32'h00000000;
assign filter_banks_5[58] = 32'h00000000;
assign filter_banks_5[59] = 32'h00000000;
assign filter_banks_5[60] = 32'h00000000;
assign filter_banks_5[61] = 32'h00000000;
assign filter_banks_5[62] = 32'h00000000;
assign filter_banks_5[63] = 32'h00000000;
assign filter_banks_5[64] = 32'h00000000;
assign filter_banks_5[65] = 32'h00000000;
assign filter_banks_5[66] = 32'h00000000;
assign filter_banks_5[67] = 32'h00000000;
assign filter_banks_5[68] = 32'h00000000;
assign filter_banks_5[69] = 32'h00000000;
assign filter_banks_5[70] = 32'h00000000;
assign filter_banks_5[71] = 32'h00000000;
assign filter_banks_5[72] = 32'h00000000;
assign filter_banks_5[73] = 32'h00000000;
assign filter_banks_5[74] = 32'h00000000;
assign filter_banks_5[75] = 32'h00000000;
assign filter_banks_5[76] = 32'h00000000;
assign filter_banks_5[77] = 32'h00000000;
assign filter_banks_5[78] = 32'h00000000;
assign filter_banks_5[79] = 32'h00000000;
assign filter_banks_5[80] = 32'h00000000;
assign filter_banks_5[81] = 32'h00000000;
assign filter_banks_5[82] = 32'h00000000;
assign filter_banks_5[83] = 32'h00000000;
assign filter_banks_5[84] = 32'h00000000;
assign filter_banks_5[85] = 32'h00000000;
assign filter_banks_5[86] = 32'h00000000;
assign filter_banks_5[87] = 32'h00000000;
assign filter_banks_5[88] = 32'h00000000;
assign filter_banks_5[89] = 32'h00000000;
assign filter_banks_5[90] = 32'h00000000;
assign filter_banks_5[91] = 32'h00000000;
assign filter_banks_5[92] = 32'h00000000;
assign filter_banks_5[93] = 32'h00000000;
assign filter_banks_5[94] = 32'h00000000;
assign filter_banks_5[95] = 32'h00000000;
assign filter_banks_5[96] = 32'h00000000;
assign filter_banks_5[97] = 32'h00000000;
assign filter_banks_5[98] = 32'h00000000;
assign filter_banks_5[99] = 32'h00000000;
assign filter_banks_5[100] = 32'h00000000;
assign filter_banks_5[101] = 32'h00000000;
assign filter_banks_5[102] = 32'h00000000;
assign filter_banks_5[103] = 32'h00000000;
assign filter_banks_5[104] = 32'h00000000;
assign filter_banks_5[105] = 32'h00000000;
assign filter_banks_5[106] = 32'h00000000;
assign filter_banks_5[107] = 32'h00000000;
assign filter_banks_5[108] = 32'h00000000;
assign filter_banks_5[109] = 32'h00000000;
assign filter_banks_5[110] = 32'h00000000;
assign filter_banks_5[111] = 32'h00000000;
assign filter_banks_5[112] = 32'h00000000;
assign filter_banks_5[113] = 32'h00000000;
assign filter_banks_5[114] = 32'h00000000;
assign filter_banks_5[115] = 32'h00000000;
assign filter_banks_5[116] = 32'h00000000;
assign filter_banks_5[117] = 32'h00000000;
assign filter_banks_5[118] = 32'h00000000;
assign filter_banks_5[119] = 32'h00000000;
assign filter_banks_5[120] = 32'h00000000;
assign filter_banks_5[121] = 32'h00000000;
assign filter_banks_5[122] = 32'h00000000;
assign filter_banks_5[123] = 32'h00000000;
assign filter_banks_5[124] = 32'h00000000;
assign filter_banks_5[125] = 32'h00000000;
assign filter_banks_5[126] = 32'h00000000;
assign filter_banks_5[127] = 32'h00000000;
assign filter_banks_5[128] = 32'h00000000;
assign filter_banks_5[129] = 32'h00000000;
assign filter_banks_5[130] = 32'h00000000;
assign filter_banks_5[131] = 32'h00000000;
assign filter_banks_5[132] = 32'h00000000;
assign filter_banks_5[133] = 32'h00000000;
assign filter_banks_5[134] = 32'h00000000;
assign filter_banks_5[135] = 32'h00000000;
assign filter_banks_5[136] = 32'h00000000;
assign filter_banks_5[137] = 32'h00000000;
assign filter_banks_5[138] = 32'h00000000;
assign filter_banks_5[139] = 32'h00000000;
assign filter_banks_5[140] = 32'h00000000;
assign filter_banks_5[141] = 32'h00000000;
assign filter_banks_5[142] = 32'h00000000;
assign filter_banks_5[143] = 32'h00000000;
assign filter_banks_5[144] = 32'h00000000;
assign filter_banks_5[145] = 32'h00000000;
assign filter_banks_5[146] = 32'h00000000;
assign filter_banks_5[147] = 32'h00000000;
assign filter_banks_5[148] = 32'h00000000;
assign filter_banks_5[149] = 32'h00000000;
assign filter_banks_5[150] = 32'h00000000;
assign filter_banks_5[151] = 32'h00000000;
assign filter_banks_5[152] = 32'h00000000;
assign filter_banks_5[153] = 32'h00000000;
assign filter_banks_5[154] = 32'h00000000;
assign filter_banks_5[155] = 32'h00000000;
assign filter_banks_5[156] = 32'h00000000;
assign filter_banks_5[157] = 32'h00000000;
assign filter_banks_5[158] = 32'h00000000;
assign filter_banks_5[159] = 32'h00000000;
assign filter_banks_5[160] = 32'h00000000;
assign filter_banks_5[161] = 32'h00000000;
assign filter_banks_5[162] = 32'h00000000;
assign filter_banks_5[163] = 32'h00000000;
assign filter_banks_5[164] = 32'h00000000;
assign filter_banks_5[165] = 32'h00000000;
assign filter_banks_5[166] = 32'h00000000;
assign filter_banks_5[167] = 32'h00000000;
assign filter_banks_5[168] = 32'h00000000;
assign filter_banks_5[169] = 32'h00000000;
assign filter_banks_5[170] = 32'h00000000;
assign filter_banks_5[171] = 32'h00000000;
assign filter_banks_5[172] = 32'h00000000;
assign filter_banks_5[173] = 32'h00000000;
assign filter_banks_5[174] = 32'h00000000;
assign filter_banks_5[175] = 32'h00000000;
assign filter_banks_5[176] = 32'h00000000;
assign filter_banks_5[177] = 32'h00000000;
assign filter_banks_5[178] = 32'h00000000;
assign filter_banks_5[179] = 32'h00000000;
assign filter_banks_5[180] = 32'h00000000;
assign filter_banks_5[181] = 32'h00000000;
assign filter_banks_5[182] = 32'h00000000;
assign filter_banks_5[183] = 32'h00000000;
assign filter_banks_5[184] = 32'h00000000;
assign filter_banks_5[185] = 32'h00000000;
assign filter_banks_5[186] = 32'h00000000;
assign filter_banks_5[187] = 32'h00000000;
assign filter_banks_5[188] = 32'h00000000;
assign filter_banks_5[189] = 32'h00000000;
assign filter_banks_5[190] = 32'h00000000;
assign filter_banks_5[191] = 32'h00000000;
assign filter_banks_5[192] = 32'h00000000;
assign filter_banks_5[193] = 32'h00000000;
assign filter_banks_5[194] = 32'h00000000;
assign filter_banks_5[195] = 32'h00000000;
assign filter_banks_5[196] = 32'h00000000;
assign filter_banks_5[197] = 32'h00000000;
assign filter_banks_5[198] = 32'h00000000;
assign filter_banks_5[199] = 32'h00000000;
assign filter_banks_5[200] = 32'h00000000;
assign filter_banks_5[201] = 32'h00000000;
assign filter_banks_5[202] = 32'h00000000;
assign filter_banks_5[203] = 32'h00000000;
assign filter_banks_5[204] = 32'h00000000;
assign filter_banks_5[205] = 32'h00000000;
assign filter_banks_5[206] = 32'h00000000;
assign filter_banks_5[207] = 32'h00000000;
assign filter_banks_5[208] = 32'h00000000;
assign filter_banks_5[209] = 32'h00000000;
assign filter_banks_5[210] = 32'h00000000;
assign filter_banks_5[211] = 32'h00000000;
assign filter_banks_5[212] = 32'h00000000;
assign filter_banks_5[213] = 32'h00000000;
assign filter_banks_5[214] = 32'h00000000;
assign filter_banks_5[215] = 32'h00000000;
assign filter_banks_5[216] = 32'h00000000;
assign filter_banks_5[217] = 32'h00000000;
assign filter_banks_5[218] = 32'h00000000;
assign filter_banks_5[219] = 32'h00000000;
assign filter_banks_5[220] = 32'h00000000;
assign filter_banks_5[221] = 32'h00000000;
assign filter_banks_5[222] = 32'h00000000;
assign filter_banks_5[223] = 32'h00000000;
assign filter_banks_5[224] = 32'h00000000;
assign filter_banks_5[225] = 32'h00000000;
assign filter_banks_5[226] = 32'h00000000;
assign filter_banks_5[227] = 32'h00000000;
assign filter_banks_5[228] = 32'h00000000;
assign filter_banks_5[229] = 32'h00000000;
assign filter_banks_5[230] = 32'h00000000;
assign filter_banks_5[231] = 32'h00000000;
assign filter_banks_5[232] = 32'h00000000;
assign filter_banks_5[233] = 32'h00000000;
assign filter_banks_5[234] = 32'h00000000;
assign filter_banks_5[235] = 32'h00000000;
assign filter_banks_5[236] = 32'h00000000;
assign filter_banks_5[237] = 32'h00000000;
assign filter_banks_5[238] = 32'h00000000;
assign filter_banks_5[239] = 32'h00000000;
assign filter_banks_5[240] = 32'h00000000;
assign filter_banks_5[241] = 32'h00000000;
assign filter_banks_5[242] = 32'h00000000;
assign filter_banks_5[243] = 32'h00000000;
assign filter_banks_5[244] = 32'h00000000;
assign filter_banks_5[245] = 32'h00000000;
assign filter_banks_5[246] = 32'h00000000;
assign filter_banks_5[247] = 32'h00000000;
assign filter_banks_5[248] = 32'h00000000;
assign filter_banks_5[249] = 32'h00000000;
assign filter_banks_5[250] = 32'h00000000;
assign filter_banks_5[251] = 32'h00000000;
assign filter_banks_5[252] = 32'h00000000;
assign filter_banks_5[253] = 32'h00000000;
assign filter_banks_5[254] = 32'h00000000;
assign filter_banks_5[255] = 32'h00000000;
assign filter_banks_5[256] = 32'h00000000;
assign filter_banks_6[0] = 32'h00000000;
assign filter_banks_6[1] = 32'h00000000;
assign filter_banks_6[2] = 32'h00000000;
assign filter_banks_6[3] = 32'h00000000;
assign filter_banks_6[4] = 32'h00000000;
assign filter_banks_6[5] = 32'h00000000;
assign filter_banks_6[6] = 32'h00000000;
assign filter_banks_6[7] = 32'h00000000;
assign filter_banks_6[8] = 32'h00000000;
assign filter_banks_6[9] = 32'h00000000;
assign filter_banks_6[10] = 32'h00000000;
assign filter_banks_6[11] = 32'h00000000;
assign filter_banks_6[12] = 32'h00000000;
assign filter_banks_6[13] = 32'h00000000;
assign filter_banks_6[14] = 32'h3eaaaaab;
assign filter_banks_6[15] = 32'h3f2aaaab;
assign filter_banks_6[16] = 32'h3f800000;
assign filter_banks_6[17] = 32'h3f400000;
assign filter_banks_6[18] = 32'h3f000000;
assign filter_banks_6[19] = 32'h3e800000;
assign filter_banks_6[20] = 32'h00000000;
assign filter_banks_6[21] = 32'h00000000;
assign filter_banks_6[22] = 32'h00000000;
assign filter_banks_6[23] = 32'h00000000;
assign filter_banks_6[24] = 32'h00000000;
assign filter_banks_6[25] = 32'h00000000;
assign filter_banks_6[26] = 32'h00000000;
assign filter_banks_6[27] = 32'h00000000;
assign filter_banks_6[28] = 32'h00000000;
assign filter_banks_6[29] = 32'h00000000;
assign filter_banks_6[30] = 32'h00000000;
assign filter_banks_6[31] = 32'h00000000;
assign filter_banks_6[32] = 32'h00000000;
assign filter_banks_6[33] = 32'h00000000;
assign filter_banks_6[34] = 32'h00000000;
assign filter_banks_6[35] = 32'h00000000;
assign filter_banks_6[36] = 32'h00000000;
assign filter_banks_6[37] = 32'h00000000;
assign filter_banks_6[38] = 32'h00000000;
assign filter_banks_6[39] = 32'h00000000;
assign filter_banks_6[40] = 32'h00000000;
assign filter_banks_6[41] = 32'h00000000;
assign filter_banks_6[42] = 32'h00000000;
assign filter_banks_6[43] = 32'h00000000;
assign filter_banks_6[44] = 32'h00000000;
assign filter_banks_6[45] = 32'h00000000;
assign filter_banks_6[46] = 32'h00000000;
assign filter_banks_6[47] = 32'h00000000;
assign filter_banks_6[48] = 32'h00000000;
assign filter_banks_6[49] = 32'h00000000;
assign filter_banks_6[50] = 32'h00000000;
assign filter_banks_6[51] = 32'h00000000;
assign filter_banks_6[52] = 32'h00000000;
assign filter_banks_6[53] = 32'h00000000;
assign filter_banks_6[54] = 32'h00000000;
assign filter_banks_6[55] = 32'h00000000;
assign filter_banks_6[56] = 32'h00000000;
assign filter_banks_6[57] = 32'h00000000;
assign filter_banks_6[58] = 32'h00000000;
assign filter_banks_6[59] = 32'h00000000;
assign filter_banks_6[60] = 32'h00000000;
assign filter_banks_6[61] = 32'h00000000;
assign filter_banks_6[62] = 32'h00000000;
assign filter_banks_6[63] = 32'h00000000;
assign filter_banks_6[64] = 32'h00000000;
assign filter_banks_6[65] = 32'h00000000;
assign filter_banks_6[66] = 32'h00000000;
assign filter_banks_6[67] = 32'h00000000;
assign filter_banks_6[68] = 32'h00000000;
assign filter_banks_6[69] = 32'h00000000;
assign filter_banks_6[70] = 32'h00000000;
assign filter_banks_6[71] = 32'h00000000;
assign filter_banks_6[72] = 32'h00000000;
assign filter_banks_6[73] = 32'h00000000;
assign filter_banks_6[74] = 32'h00000000;
assign filter_banks_6[75] = 32'h00000000;
assign filter_banks_6[76] = 32'h00000000;
assign filter_banks_6[77] = 32'h00000000;
assign filter_banks_6[78] = 32'h00000000;
assign filter_banks_6[79] = 32'h00000000;
assign filter_banks_6[80] = 32'h00000000;
assign filter_banks_6[81] = 32'h00000000;
assign filter_banks_6[82] = 32'h00000000;
assign filter_banks_6[83] = 32'h00000000;
assign filter_banks_6[84] = 32'h00000000;
assign filter_banks_6[85] = 32'h00000000;
assign filter_banks_6[86] = 32'h00000000;
assign filter_banks_6[87] = 32'h00000000;
assign filter_banks_6[88] = 32'h00000000;
assign filter_banks_6[89] = 32'h00000000;
assign filter_banks_6[90] = 32'h00000000;
assign filter_banks_6[91] = 32'h00000000;
assign filter_banks_6[92] = 32'h00000000;
assign filter_banks_6[93] = 32'h00000000;
assign filter_banks_6[94] = 32'h00000000;
assign filter_banks_6[95] = 32'h00000000;
assign filter_banks_6[96] = 32'h00000000;
assign filter_banks_6[97] = 32'h00000000;
assign filter_banks_6[98] = 32'h00000000;
assign filter_banks_6[99] = 32'h00000000;
assign filter_banks_6[100] = 32'h00000000;
assign filter_banks_6[101] = 32'h00000000;
assign filter_banks_6[102] = 32'h00000000;
assign filter_banks_6[103] = 32'h00000000;
assign filter_banks_6[104] = 32'h00000000;
assign filter_banks_6[105] = 32'h00000000;
assign filter_banks_6[106] = 32'h00000000;
assign filter_banks_6[107] = 32'h00000000;
assign filter_banks_6[108] = 32'h00000000;
assign filter_banks_6[109] = 32'h00000000;
assign filter_banks_6[110] = 32'h00000000;
assign filter_banks_6[111] = 32'h00000000;
assign filter_banks_6[112] = 32'h00000000;
assign filter_banks_6[113] = 32'h00000000;
assign filter_banks_6[114] = 32'h00000000;
assign filter_banks_6[115] = 32'h00000000;
assign filter_banks_6[116] = 32'h00000000;
assign filter_banks_6[117] = 32'h00000000;
assign filter_banks_6[118] = 32'h00000000;
assign filter_banks_6[119] = 32'h00000000;
assign filter_banks_6[120] = 32'h00000000;
assign filter_banks_6[121] = 32'h00000000;
assign filter_banks_6[122] = 32'h00000000;
assign filter_banks_6[123] = 32'h00000000;
assign filter_banks_6[124] = 32'h00000000;
assign filter_banks_6[125] = 32'h00000000;
assign filter_banks_6[126] = 32'h00000000;
assign filter_banks_6[127] = 32'h00000000;
assign filter_banks_6[128] = 32'h00000000;
assign filter_banks_6[129] = 32'h00000000;
assign filter_banks_6[130] = 32'h00000000;
assign filter_banks_6[131] = 32'h00000000;
assign filter_banks_6[132] = 32'h00000000;
assign filter_banks_6[133] = 32'h00000000;
assign filter_banks_6[134] = 32'h00000000;
assign filter_banks_6[135] = 32'h00000000;
assign filter_banks_6[136] = 32'h00000000;
assign filter_banks_6[137] = 32'h00000000;
assign filter_banks_6[138] = 32'h00000000;
assign filter_banks_6[139] = 32'h00000000;
assign filter_banks_6[140] = 32'h00000000;
assign filter_banks_6[141] = 32'h00000000;
assign filter_banks_6[142] = 32'h00000000;
assign filter_banks_6[143] = 32'h00000000;
assign filter_banks_6[144] = 32'h00000000;
assign filter_banks_6[145] = 32'h00000000;
assign filter_banks_6[146] = 32'h00000000;
assign filter_banks_6[147] = 32'h00000000;
assign filter_banks_6[148] = 32'h00000000;
assign filter_banks_6[149] = 32'h00000000;
assign filter_banks_6[150] = 32'h00000000;
assign filter_banks_6[151] = 32'h00000000;
assign filter_banks_6[152] = 32'h00000000;
assign filter_banks_6[153] = 32'h00000000;
assign filter_banks_6[154] = 32'h00000000;
assign filter_banks_6[155] = 32'h00000000;
assign filter_banks_6[156] = 32'h00000000;
assign filter_banks_6[157] = 32'h00000000;
assign filter_banks_6[158] = 32'h00000000;
assign filter_banks_6[159] = 32'h00000000;
assign filter_banks_6[160] = 32'h00000000;
assign filter_banks_6[161] = 32'h00000000;
assign filter_banks_6[162] = 32'h00000000;
assign filter_banks_6[163] = 32'h00000000;
assign filter_banks_6[164] = 32'h00000000;
assign filter_banks_6[165] = 32'h00000000;
assign filter_banks_6[166] = 32'h00000000;
assign filter_banks_6[167] = 32'h00000000;
assign filter_banks_6[168] = 32'h00000000;
assign filter_banks_6[169] = 32'h00000000;
assign filter_banks_6[170] = 32'h00000000;
assign filter_banks_6[171] = 32'h00000000;
assign filter_banks_6[172] = 32'h00000000;
assign filter_banks_6[173] = 32'h00000000;
assign filter_banks_6[174] = 32'h00000000;
assign filter_banks_6[175] = 32'h00000000;
assign filter_banks_6[176] = 32'h00000000;
assign filter_banks_6[177] = 32'h00000000;
assign filter_banks_6[178] = 32'h00000000;
assign filter_banks_6[179] = 32'h00000000;
assign filter_banks_6[180] = 32'h00000000;
assign filter_banks_6[181] = 32'h00000000;
assign filter_banks_6[182] = 32'h00000000;
assign filter_banks_6[183] = 32'h00000000;
assign filter_banks_6[184] = 32'h00000000;
assign filter_banks_6[185] = 32'h00000000;
assign filter_banks_6[186] = 32'h00000000;
assign filter_banks_6[187] = 32'h00000000;
assign filter_banks_6[188] = 32'h00000000;
assign filter_banks_6[189] = 32'h00000000;
assign filter_banks_6[190] = 32'h00000000;
assign filter_banks_6[191] = 32'h00000000;
assign filter_banks_6[192] = 32'h00000000;
assign filter_banks_6[193] = 32'h00000000;
assign filter_banks_6[194] = 32'h00000000;
assign filter_banks_6[195] = 32'h00000000;
assign filter_banks_6[196] = 32'h00000000;
assign filter_banks_6[197] = 32'h00000000;
assign filter_banks_6[198] = 32'h00000000;
assign filter_banks_6[199] = 32'h00000000;
assign filter_banks_6[200] = 32'h00000000;
assign filter_banks_6[201] = 32'h00000000;
assign filter_banks_6[202] = 32'h00000000;
assign filter_banks_6[203] = 32'h00000000;
assign filter_banks_6[204] = 32'h00000000;
assign filter_banks_6[205] = 32'h00000000;
assign filter_banks_6[206] = 32'h00000000;
assign filter_banks_6[207] = 32'h00000000;
assign filter_banks_6[208] = 32'h00000000;
assign filter_banks_6[209] = 32'h00000000;
assign filter_banks_6[210] = 32'h00000000;
assign filter_banks_6[211] = 32'h00000000;
assign filter_banks_6[212] = 32'h00000000;
assign filter_banks_6[213] = 32'h00000000;
assign filter_banks_6[214] = 32'h00000000;
assign filter_banks_6[215] = 32'h00000000;
assign filter_banks_6[216] = 32'h00000000;
assign filter_banks_6[217] = 32'h00000000;
assign filter_banks_6[218] = 32'h00000000;
assign filter_banks_6[219] = 32'h00000000;
assign filter_banks_6[220] = 32'h00000000;
assign filter_banks_6[221] = 32'h00000000;
assign filter_banks_6[222] = 32'h00000000;
assign filter_banks_6[223] = 32'h00000000;
assign filter_banks_6[224] = 32'h00000000;
assign filter_banks_6[225] = 32'h00000000;
assign filter_banks_6[226] = 32'h00000000;
assign filter_banks_6[227] = 32'h00000000;
assign filter_banks_6[228] = 32'h00000000;
assign filter_banks_6[229] = 32'h00000000;
assign filter_banks_6[230] = 32'h00000000;
assign filter_banks_6[231] = 32'h00000000;
assign filter_banks_6[232] = 32'h00000000;
assign filter_banks_6[233] = 32'h00000000;
assign filter_banks_6[234] = 32'h00000000;
assign filter_banks_6[235] = 32'h00000000;
assign filter_banks_6[236] = 32'h00000000;
assign filter_banks_6[237] = 32'h00000000;
assign filter_banks_6[238] = 32'h00000000;
assign filter_banks_6[239] = 32'h00000000;
assign filter_banks_6[240] = 32'h00000000;
assign filter_banks_6[241] = 32'h00000000;
assign filter_banks_6[242] = 32'h00000000;
assign filter_banks_6[243] = 32'h00000000;
assign filter_banks_6[244] = 32'h00000000;
assign filter_banks_6[245] = 32'h00000000;
assign filter_banks_6[246] = 32'h00000000;
assign filter_banks_6[247] = 32'h00000000;
assign filter_banks_6[248] = 32'h00000000;
assign filter_banks_6[249] = 32'h00000000;
assign filter_banks_6[250] = 32'h00000000;
assign filter_banks_6[251] = 32'h00000000;
assign filter_banks_6[252] = 32'h00000000;
assign filter_banks_6[253] = 32'h00000000;
assign filter_banks_6[254] = 32'h00000000;
assign filter_banks_6[255] = 32'h00000000;
assign filter_banks_6[256] = 32'h00000000;
assign filter_banks_7[0] = 32'h00000000;
assign filter_banks_7[1] = 32'h00000000;
assign filter_banks_7[2] = 32'h00000000;
assign filter_banks_7[3] = 32'h00000000;
assign filter_banks_7[4] = 32'h00000000;
assign filter_banks_7[5] = 32'h00000000;
assign filter_banks_7[6] = 32'h00000000;
assign filter_banks_7[7] = 32'h00000000;
assign filter_banks_7[8] = 32'h00000000;
assign filter_banks_7[9] = 32'h00000000;
assign filter_banks_7[10] = 32'h00000000;
assign filter_banks_7[11] = 32'h00000000;
assign filter_banks_7[12] = 32'h00000000;
assign filter_banks_7[13] = 32'h00000000;
assign filter_banks_7[14] = 32'h00000000;
assign filter_banks_7[15] = 32'h00000000;
assign filter_banks_7[16] = 32'h00000000;
assign filter_banks_7[17] = 32'h3e800000;
assign filter_banks_7[18] = 32'h3f000000;
assign filter_banks_7[19] = 32'h3f400000;
assign filter_banks_7[20] = 32'h3f800000;
assign filter_banks_7[21] = 32'h3f400000;
assign filter_banks_7[22] = 32'h3f000000;
assign filter_banks_7[23] = 32'h3e800000;
assign filter_banks_7[24] = 32'h00000000;
assign filter_banks_7[25] = 32'h00000000;
assign filter_banks_7[26] = 32'h00000000;
assign filter_banks_7[27] = 32'h00000000;
assign filter_banks_7[28] = 32'h00000000;
assign filter_banks_7[29] = 32'h00000000;
assign filter_banks_7[30] = 32'h00000000;
assign filter_banks_7[31] = 32'h00000000;
assign filter_banks_7[32] = 32'h00000000;
assign filter_banks_7[33] = 32'h00000000;
assign filter_banks_7[34] = 32'h00000000;
assign filter_banks_7[35] = 32'h00000000;
assign filter_banks_7[36] = 32'h00000000;
assign filter_banks_7[37] = 32'h00000000;
assign filter_banks_7[38] = 32'h00000000;
assign filter_banks_7[39] = 32'h00000000;
assign filter_banks_7[40] = 32'h00000000;
assign filter_banks_7[41] = 32'h00000000;
assign filter_banks_7[42] = 32'h00000000;
assign filter_banks_7[43] = 32'h00000000;
assign filter_banks_7[44] = 32'h00000000;
assign filter_banks_7[45] = 32'h00000000;
assign filter_banks_7[46] = 32'h00000000;
assign filter_banks_7[47] = 32'h00000000;
assign filter_banks_7[48] = 32'h00000000;
assign filter_banks_7[49] = 32'h00000000;
assign filter_banks_7[50] = 32'h00000000;
assign filter_banks_7[51] = 32'h00000000;
assign filter_banks_7[52] = 32'h00000000;
assign filter_banks_7[53] = 32'h00000000;
assign filter_banks_7[54] = 32'h00000000;
assign filter_banks_7[55] = 32'h00000000;
assign filter_banks_7[56] = 32'h00000000;
assign filter_banks_7[57] = 32'h00000000;
assign filter_banks_7[58] = 32'h00000000;
assign filter_banks_7[59] = 32'h00000000;
assign filter_banks_7[60] = 32'h00000000;
assign filter_banks_7[61] = 32'h00000000;
assign filter_banks_7[62] = 32'h00000000;
assign filter_banks_7[63] = 32'h00000000;
assign filter_banks_7[64] = 32'h00000000;
assign filter_banks_7[65] = 32'h00000000;
assign filter_banks_7[66] = 32'h00000000;
assign filter_banks_7[67] = 32'h00000000;
assign filter_banks_7[68] = 32'h00000000;
assign filter_banks_7[69] = 32'h00000000;
assign filter_banks_7[70] = 32'h00000000;
assign filter_banks_7[71] = 32'h00000000;
assign filter_banks_7[72] = 32'h00000000;
assign filter_banks_7[73] = 32'h00000000;
assign filter_banks_7[74] = 32'h00000000;
assign filter_banks_7[75] = 32'h00000000;
assign filter_banks_7[76] = 32'h00000000;
assign filter_banks_7[77] = 32'h00000000;
assign filter_banks_7[78] = 32'h00000000;
assign filter_banks_7[79] = 32'h00000000;
assign filter_banks_7[80] = 32'h00000000;
assign filter_banks_7[81] = 32'h00000000;
assign filter_banks_7[82] = 32'h00000000;
assign filter_banks_7[83] = 32'h00000000;
assign filter_banks_7[84] = 32'h00000000;
assign filter_banks_7[85] = 32'h00000000;
assign filter_banks_7[86] = 32'h00000000;
assign filter_banks_7[87] = 32'h00000000;
assign filter_banks_7[88] = 32'h00000000;
assign filter_banks_7[89] = 32'h00000000;
assign filter_banks_7[90] = 32'h00000000;
assign filter_banks_7[91] = 32'h00000000;
assign filter_banks_7[92] = 32'h00000000;
assign filter_banks_7[93] = 32'h00000000;
assign filter_banks_7[94] = 32'h00000000;
assign filter_banks_7[95] = 32'h00000000;
assign filter_banks_7[96] = 32'h00000000;
assign filter_banks_7[97] = 32'h00000000;
assign filter_banks_7[98] = 32'h00000000;
assign filter_banks_7[99] = 32'h00000000;
assign filter_banks_7[100] = 32'h00000000;
assign filter_banks_7[101] = 32'h00000000;
assign filter_banks_7[102] = 32'h00000000;
assign filter_banks_7[103] = 32'h00000000;
assign filter_banks_7[104] = 32'h00000000;
assign filter_banks_7[105] = 32'h00000000;
assign filter_banks_7[106] = 32'h00000000;
assign filter_banks_7[107] = 32'h00000000;
assign filter_banks_7[108] = 32'h00000000;
assign filter_banks_7[109] = 32'h00000000;
assign filter_banks_7[110] = 32'h00000000;
assign filter_banks_7[111] = 32'h00000000;
assign filter_banks_7[112] = 32'h00000000;
assign filter_banks_7[113] = 32'h00000000;
assign filter_banks_7[114] = 32'h00000000;
assign filter_banks_7[115] = 32'h00000000;
assign filter_banks_7[116] = 32'h00000000;
assign filter_banks_7[117] = 32'h00000000;
assign filter_banks_7[118] = 32'h00000000;
assign filter_banks_7[119] = 32'h00000000;
assign filter_banks_7[120] = 32'h00000000;
assign filter_banks_7[121] = 32'h00000000;
assign filter_banks_7[122] = 32'h00000000;
assign filter_banks_7[123] = 32'h00000000;
assign filter_banks_7[124] = 32'h00000000;
assign filter_banks_7[125] = 32'h00000000;
assign filter_banks_7[126] = 32'h00000000;
assign filter_banks_7[127] = 32'h00000000;
assign filter_banks_7[128] = 32'h00000000;
assign filter_banks_7[129] = 32'h00000000;
assign filter_banks_7[130] = 32'h00000000;
assign filter_banks_7[131] = 32'h00000000;
assign filter_banks_7[132] = 32'h00000000;
assign filter_banks_7[133] = 32'h00000000;
assign filter_banks_7[134] = 32'h00000000;
assign filter_banks_7[135] = 32'h00000000;
assign filter_banks_7[136] = 32'h00000000;
assign filter_banks_7[137] = 32'h00000000;
assign filter_banks_7[138] = 32'h00000000;
assign filter_banks_7[139] = 32'h00000000;
assign filter_banks_7[140] = 32'h00000000;
assign filter_banks_7[141] = 32'h00000000;
assign filter_banks_7[142] = 32'h00000000;
assign filter_banks_7[143] = 32'h00000000;
assign filter_banks_7[144] = 32'h00000000;
assign filter_banks_7[145] = 32'h00000000;
assign filter_banks_7[146] = 32'h00000000;
assign filter_banks_7[147] = 32'h00000000;
assign filter_banks_7[148] = 32'h00000000;
assign filter_banks_7[149] = 32'h00000000;
assign filter_banks_7[150] = 32'h00000000;
assign filter_banks_7[151] = 32'h00000000;
assign filter_banks_7[152] = 32'h00000000;
assign filter_banks_7[153] = 32'h00000000;
assign filter_banks_7[154] = 32'h00000000;
assign filter_banks_7[155] = 32'h00000000;
assign filter_banks_7[156] = 32'h00000000;
assign filter_banks_7[157] = 32'h00000000;
assign filter_banks_7[158] = 32'h00000000;
assign filter_banks_7[159] = 32'h00000000;
assign filter_banks_7[160] = 32'h00000000;
assign filter_banks_7[161] = 32'h00000000;
assign filter_banks_7[162] = 32'h00000000;
assign filter_banks_7[163] = 32'h00000000;
assign filter_banks_7[164] = 32'h00000000;
assign filter_banks_7[165] = 32'h00000000;
assign filter_banks_7[166] = 32'h00000000;
assign filter_banks_7[167] = 32'h00000000;
assign filter_banks_7[168] = 32'h00000000;
assign filter_banks_7[169] = 32'h00000000;
assign filter_banks_7[170] = 32'h00000000;
assign filter_banks_7[171] = 32'h00000000;
assign filter_banks_7[172] = 32'h00000000;
assign filter_banks_7[173] = 32'h00000000;
assign filter_banks_7[174] = 32'h00000000;
assign filter_banks_7[175] = 32'h00000000;
assign filter_banks_7[176] = 32'h00000000;
assign filter_banks_7[177] = 32'h00000000;
assign filter_banks_7[178] = 32'h00000000;
assign filter_banks_7[179] = 32'h00000000;
assign filter_banks_7[180] = 32'h00000000;
assign filter_banks_7[181] = 32'h00000000;
assign filter_banks_7[182] = 32'h00000000;
assign filter_banks_7[183] = 32'h00000000;
assign filter_banks_7[184] = 32'h00000000;
assign filter_banks_7[185] = 32'h00000000;
assign filter_banks_7[186] = 32'h00000000;
assign filter_banks_7[187] = 32'h00000000;
assign filter_banks_7[188] = 32'h00000000;
assign filter_banks_7[189] = 32'h00000000;
assign filter_banks_7[190] = 32'h00000000;
assign filter_banks_7[191] = 32'h00000000;
assign filter_banks_7[192] = 32'h00000000;
assign filter_banks_7[193] = 32'h00000000;
assign filter_banks_7[194] = 32'h00000000;
assign filter_banks_7[195] = 32'h00000000;
assign filter_banks_7[196] = 32'h00000000;
assign filter_banks_7[197] = 32'h00000000;
assign filter_banks_7[198] = 32'h00000000;
assign filter_banks_7[199] = 32'h00000000;
assign filter_banks_7[200] = 32'h00000000;
assign filter_banks_7[201] = 32'h00000000;
assign filter_banks_7[202] = 32'h00000000;
assign filter_banks_7[203] = 32'h00000000;
assign filter_banks_7[204] = 32'h00000000;
assign filter_banks_7[205] = 32'h00000000;
assign filter_banks_7[206] = 32'h00000000;
assign filter_banks_7[207] = 32'h00000000;
assign filter_banks_7[208] = 32'h00000000;
assign filter_banks_7[209] = 32'h00000000;
assign filter_banks_7[210] = 32'h00000000;
assign filter_banks_7[211] = 32'h00000000;
assign filter_banks_7[212] = 32'h00000000;
assign filter_banks_7[213] = 32'h00000000;
assign filter_banks_7[214] = 32'h00000000;
assign filter_banks_7[215] = 32'h00000000;
assign filter_banks_7[216] = 32'h00000000;
assign filter_banks_7[217] = 32'h00000000;
assign filter_banks_7[218] = 32'h00000000;
assign filter_banks_7[219] = 32'h00000000;
assign filter_banks_7[220] = 32'h00000000;
assign filter_banks_7[221] = 32'h00000000;
assign filter_banks_7[222] = 32'h00000000;
assign filter_banks_7[223] = 32'h00000000;
assign filter_banks_7[224] = 32'h00000000;
assign filter_banks_7[225] = 32'h00000000;
assign filter_banks_7[226] = 32'h00000000;
assign filter_banks_7[227] = 32'h00000000;
assign filter_banks_7[228] = 32'h00000000;
assign filter_banks_7[229] = 32'h00000000;
assign filter_banks_7[230] = 32'h00000000;
assign filter_banks_7[231] = 32'h00000000;
assign filter_banks_7[232] = 32'h00000000;
assign filter_banks_7[233] = 32'h00000000;
assign filter_banks_7[234] = 32'h00000000;
assign filter_banks_7[235] = 32'h00000000;
assign filter_banks_7[236] = 32'h00000000;
assign filter_banks_7[237] = 32'h00000000;
assign filter_banks_7[238] = 32'h00000000;
assign filter_banks_7[239] = 32'h00000000;
assign filter_banks_7[240] = 32'h00000000;
assign filter_banks_7[241] = 32'h00000000;
assign filter_banks_7[242] = 32'h00000000;
assign filter_banks_7[243] = 32'h00000000;
assign filter_banks_7[244] = 32'h00000000;
assign filter_banks_7[245] = 32'h00000000;
assign filter_banks_7[246] = 32'h00000000;
assign filter_banks_7[247] = 32'h00000000;
assign filter_banks_7[248] = 32'h00000000;
assign filter_banks_7[249] = 32'h00000000;
assign filter_banks_7[250] = 32'h00000000;
assign filter_banks_7[251] = 32'h00000000;
assign filter_banks_7[252] = 32'h00000000;
assign filter_banks_7[253] = 32'h00000000;
assign filter_banks_7[254] = 32'h00000000;
assign filter_banks_7[255] = 32'h00000000;
assign filter_banks_7[256] = 32'h00000000;
assign filter_banks_8[0] = 32'h00000000;
assign filter_banks_8[1] = 32'h00000000;
assign filter_banks_8[2] = 32'h00000000;
assign filter_banks_8[3] = 32'h00000000;
assign filter_banks_8[4] = 32'h00000000;
assign filter_banks_8[5] = 32'h00000000;
assign filter_banks_8[6] = 32'h00000000;
assign filter_banks_8[7] = 32'h00000000;
assign filter_banks_8[8] = 32'h00000000;
assign filter_banks_8[9] = 32'h00000000;
assign filter_banks_8[10] = 32'h00000000;
assign filter_banks_8[11] = 32'h00000000;
assign filter_banks_8[12] = 32'h00000000;
assign filter_banks_8[13] = 32'h00000000;
assign filter_banks_8[14] = 32'h00000000;
assign filter_banks_8[15] = 32'h00000000;
assign filter_banks_8[16] = 32'h00000000;
assign filter_banks_8[17] = 32'h00000000;
assign filter_banks_8[18] = 32'h00000000;
assign filter_banks_8[19] = 32'h00000000;
assign filter_banks_8[20] = 32'h00000000;
assign filter_banks_8[21] = 32'h3e800000;
assign filter_banks_8[22] = 32'h3f000000;
assign filter_banks_8[23] = 32'h3f400000;
assign filter_banks_8[24] = 32'h3f800000;
assign filter_banks_8[25] = 32'h3f4ccccd;
assign filter_banks_8[26] = 32'h3f19999a;
assign filter_banks_8[27] = 32'h3ecccccd;
assign filter_banks_8[28] = 32'h3e4ccccd;
assign filter_banks_8[29] = 32'h00000000;
assign filter_banks_8[30] = 32'h00000000;
assign filter_banks_8[31] = 32'h00000000;
assign filter_banks_8[32] = 32'h00000000;
assign filter_banks_8[33] = 32'h00000000;
assign filter_banks_8[34] = 32'h00000000;
assign filter_banks_8[35] = 32'h00000000;
assign filter_banks_8[36] = 32'h00000000;
assign filter_banks_8[37] = 32'h00000000;
assign filter_banks_8[38] = 32'h00000000;
assign filter_banks_8[39] = 32'h00000000;
assign filter_banks_8[40] = 32'h00000000;
assign filter_banks_8[41] = 32'h00000000;
assign filter_banks_8[42] = 32'h00000000;
assign filter_banks_8[43] = 32'h00000000;
assign filter_banks_8[44] = 32'h00000000;
assign filter_banks_8[45] = 32'h00000000;
assign filter_banks_8[46] = 32'h00000000;
assign filter_banks_8[47] = 32'h00000000;
assign filter_banks_8[48] = 32'h00000000;
assign filter_banks_8[49] = 32'h00000000;
assign filter_banks_8[50] = 32'h00000000;
assign filter_banks_8[51] = 32'h00000000;
assign filter_banks_8[52] = 32'h00000000;
assign filter_banks_8[53] = 32'h00000000;
assign filter_banks_8[54] = 32'h00000000;
assign filter_banks_8[55] = 32'h00000000;
assign filter_banks_8[56] = 32'h00000000;
assign filter_banks_8[57] = 32'h00000000;
assign filter_banks_8[58] = 32'h00000000;
assign filter_banks_8[59] = 32'h00000000;
assign filter_banks_8[60] = 32'h00000000;
assign filter_banks_8[61] = 32'h00000000;
assign filter_banks_8[62] = 32'h00000000;
assign filter_banks_8[63] = 32'h00000000;
assign filter_banks_8[64] = 32'h00000000;
assign filter_banks_8[65] = 32'h00000000;
assign filter_banks_8[66] = 32'h00000000;
assign filter_banks_8[67] = 32'h00000000;
assign filter_banks_8[68] = 32'h00000000;
assign filter_banks_8[69] = 32'h00000000;
assign filter_banks_8[70] = 32'h00000000;
assign filter_banks_8[71] = 32'h00000000;
assign filter_banks_8[72] = 32'h00000000;
assign filter_banks_8[73] = 32'h00000000;
assign filter_banks_8[74] = 32'h00000000;
assign filter_banks_8[75] = 32'h00000000;
assign filter_banks_8[76] = 32'h00000000;
assign filter_banks_8[77] = 32'h00000000;
assign filter_banks_8[78] = 32'h00000000;
assign filter_banks_8[79] = 32'h00000000;
assign filter_banks_8[80] = 32'h00000000;
assign filter_banks_8[81] = 32'h00000000;
assign filter_banks_8[82] = 32'h00000000;
assign filter_banks_8[83] = 32'h00000000;
assign filter_banks_8[84] = 32'h00000000;
assign filter_banks_8[85] = 32'h00000000;
assign filter_banks_8[86] = 32'h00000000;
assign filter_banks_8[87] = 32'h00000000;
assign filter_banks_8[88] = 32'h00000000;
assign filter_banks_8[89] = 32'h00000000;
assign filter_banks_8[90] = 32'h00000000;
assign filter_banks_8[91] = 32'h00000000;
assign filter_banks_8[92] = 32'h00000000;
assign filter_banks_8[93] = 32'h00000000;
assign filter_banks_8[94] = 32'h00000000;
assign filter_banks_8[95] = 32'h00000000;
assign filter_banks_8[96] = 32'h00000000;
assign filter_banks_8[97] = 32'h00000000;
assign filter_banks_8[98] = 32'h00000000;
assign filter_banks_8[99] = 32'h00000000;
assign filter_banks_8[100] = 32'h00000000;
assign filter_banks_8[101] = 32'h00000000;
assign filter_banks_8[102] = 32'h00000000;
assign filter_banks_8[103] = 32'h00000000;
assign filter_banks_8[104] = 32'h00000000;
assign filter_banks_8[105] = 32'h00000000;
assign filter_banks_8[106] = 32'h00000000;
assign filter_banks_8[107] = 32'h00000000;
assign filter_banks_8[108] = 32'h00000000;
assign filter_banks_8[109] = 32'h00000000;
assign filter_banks_8[110] = 32'h00000000;
assign filter_banks_8[111] = 32'h00000000;
assign filter_banks_8[112] = 32'h00000000;
assign filter_banks_8[113] = 32'h00000000;
assign filter_banks_8[114] = 32'h00000000;
assign filter_banks_8[115] = 32'h00000000;
assign filter_banks_8[116] = 32'h00000000;
assign filter_banks_8[117] = 32'h00000000;
assign filter_banks_8[118] = 32'h00000000;
assign filter_banks_8[119] = 32'h00000000;
assign filter_banks_8[120] = 32'h00000000;
assign filter_banks_8[121] = 32'h00000000;
assign filter_banks_8[122] = 32'h00000000;
assign filter_banks_8[123] = 32'h00000000;
assign filter_banks_8[124] = 32'h00000000;
assign filter_banks_8[125] = 32'h00000000;
assign filter_banks_8[126] = 32'h00000000;
assign filter_banks_8[127] = 32'h00000000;
assign filter_banks_8[128] = 32'h00000000;
assign filter_banks_8[129] = 32'h00000000;
assign filter_banks_8[130] = 32'h00000000;
assign filter_banks_8[131] = 32'h00000000;
assign filter_banks_8[132] = 32'h00000000;
assign filter_banks_8[133] = 32'h00000000;
assign filter_banks_8[134] = 32'h00000000;
assign filter_banks_8[135] = 32'h00000000;
assign filter_banks_8[136] = 32'h00000000;
assign filter_banks_8[137] = 32'h00000000;
assign filter_banks_8[138] = 32'h00000000;
assign filter_banks_8[139] = 32'h00000000;
assign filter_banks_8[140] = 32'h00000000;
assign filter_banks_8[141] = 32'h00000000;
assign filter_banks_8[142] = 32'h00000000;
assign filter_banks_8[143] = 32'h00000000;
assign filter_banks_8[144] = 32'h00000000;
assign filter_banks_8[145] = 32'h00000000;
assign filter_banks_8[146] = 32'h00000000;
assign filter_banks_8[147] = 32'h00000000;
assign filter_banks_8[148] = 32'h00000000;
assign filter_banks_8[149] = 32'h00000000;
assign filter_banks_8[150] = 32'h00000000;
assign filter_banks_8[151] = 32'h00000000;
assign filter_banks_8[152] = 32'h00000000;
assign filter_banks_8[153] = 32'h00000000;
assign filter_banks_8[154] = 32'h00000000;
assign filter_banks_8[155] = 32'h00000000;
assign filter_banks_8[156] = 32'h00000000;
assign filter_banks_8[157] = 32'h00000000;
assign filter_banks_8[158] = 32'h00000000;
assign filter_banks_8[159] = 32'h00000000;
assign filter_banks_8[160] = 32'h00000000;
assign filter_banks_8[161] = 32'h00000000;
assign filter_banks_8[162] = 32'h00000000;
assign filter_banks_8[163] = 32'h00000000;
assign filter_banks_8[164] = 32'h00000000;
assign filter_banks_8[165] = 32'h00000000;
assign filter_banks_8[166] = 32'h00000000;
assign filter_banks_8[167] = 32'h00000000;
assign filter_banks_8[168] = 32'h00000000;
assign filter_banks_8[169] = 32'h00000000;
assign filter_banks_8[170] = 32'h00000000;
assign filter_banks_8[171] = 32'h00000000;
assign filter_banks_8[172] = 32'h00000000;
assign filter_banks_8[173] = 32'h00000000;
assign filter_banks_8[174] = 32'h00000000;
assign filter_banks_8[175] = 32'h00000000;
assign filter_banks_8[176] = 32'h00000000;
assign filter_banks_8[177] = 32'h00000000;
assign filter_banks_8[178] = 32'h00000000;
assign filter_banks_8[179] = 32'h00000000;
assign filter_banks_8[180] = 32'h00000000;
assign filter_banks_8[181] = 32'h00000000;
assign filter_banks_8[182] = 32'h00000000;
assign filter_banks_8[183] = 32'h00000000;
assign filter_banks_8[184] = 32'h00000000;
assign filter_banks_8[185] = 32'h00000000;
assign filter_banks_8[186] = 32'h00000000;
assign filter_banks_8[187] = 32'h00000000;
assign filter_banks_8[188] = 32'h00000000;
assign filter_banks_8[189] = 32'h00000000;
assign filter_banks_8[190] = 32'h00000000;
assign filter_banks_8[191] = 32'h00000000;
assign filter_banks_8[192] = 32'h00000000;
assign filter_banks_8[193] = 32'h00000000;
assign filter_banks_8[194] = 32'h00000000;
assign filter_banks_8[195] = 32'h00000000;
assign filter_banks_8[196] = 32'h00000000;
assign filter_banks_8[197] = 32'h00000000;
assign filter_banks_8[198] = 32'h00000000;
assign filter_banks_8[199] = 32'h00000000;
assign filter_banks_8[200] = 32'h00000000;
assign filter_banks_8[201] = 32'h00000000;
assign filter_banks_8[202] = 32'h00000000;
assign filter_banks_8[203] = 32'h00000000;
assign filter_banks_8[204] = 32'h00000000;
assign filter_banks_8[205] = 32'h00000000;
assign filter_banks_8[206] = 32'h00000000;
assign filter_banks_8[207] = 32'h00000000;
assign filter_banks_8[208] = 32'h00000000;
assign filter_banks_8[209] = 32'h00000000;
assign filter_banks_8[210] = 32'h00000000;
assign filter_banks_8[211] = 32'h00000000;
assign filter_banks_8[212] = 32'h00000000;
assign filter_banks_8[213] = 32'h00000000;
assign filter_banks_8[214] = 32'h00000000;
assign filter_banks_8[215] = 32'h00000000;
assign filter_banks_8[216] = 32'h00000000;
assign filter_banks_8[217] = 32'h00000000;
assign filter_banks_8[218] = 32'h00000000;
assign filter_banks_8[219] = 32'h00000000;
assign filter_banks_8[220] = 32'h00000000;
assign filter_banks_8[221] = 32'h00000000;
assign filter_banks_8[222] = 32'h00000000;
assign filter_banks_8[223] = 32'h00000000;
assign filter_banks_8[224] = 32'h00000000;
assign filter_banks_8[225] = 32'h00000000;
assign filter_banks_8[226] = 32'h00000000;
assign filter_banks_8[227] = 32'h00000000;
assign filter_banks_8[228] = 32'h00000000;
assign filter_banks_8[229] = 32'h00000000;
assign filter_banks_8[230] = 32'h00000000;
assign filter_banks_8[231] = 32'h00000000;
assign filter_banks_8[232] = 32'h00000000;
assign filter_banks_8[233] = 32'h00000000;
assign filter_banks_8[234] = 32'h00000000;
assign filter_banks_8[235] = 32'h00000000;
assign filter_banks_8[236] = 32'h00000000;
assign filter_banks_8[237] = 32'h00000000;
assign filter_banks_8[238] = 32'h00000000;
assign filter_banks_8[239] = 32'h00000000;
assign filter_banks_8[240] = 32'h00000000;
assign filter_banks_8[241] = 32'h00000000;
assign filter_banks_8[242] = 32'h00000000;
assign filter_banks_8[243] = 32'h00000000;
assign filter_banks_8[244] = 32'h00000000;
assign filter_banks_8[245] = 32'h00000000;
assign filter_banks_8[246] = 32'h00000000;
assign filter_banks_8[247] = 32'h00000000;
assign filter_banks_8[248] = 32'h00000000;
assign filter_banks_8[249] = 32'h00000000;
assign filter_banks_8[250] = 32'h00000000;
assign filter_banks_8[251] = 32'h00000000;
assign filter_banks_8[252] = 32'h00000000;
assign filter_banks_8[253] = 32'h00000000;
assign filter_banks_8[254] = 32'h00000000;
assign filter_banks_8[255] = 32'h00000000;
assign filter_banks_8[256] = 32'h00000000;
assign filter_banks_9[0] = 32'h00000000;
assign filter_banks_9[1] = 32'h00000000;
assign filter_banks_9[2] = 32'h00000000;
assign filter_banks_9[3] = 32'h00000000;
assign filter_banks_9[4] = 32'h00000000;
assign filter_banks_9[5] = 32'h00000000;
assign filter_banks_9[6] = 32'h00000000;
assign filter_banks_9[7] = 32'h00000000;
assign filter_banks_9[8] = 32'h00000000;
assign filter_banks_9[9] = 32'h00000000;
assign filter_banks_9[10] = 32'h00000000;
assign filter_banks_9[11] = 32'h00000000;
assign filter_banks_9[12] = 32'h00000000;
assign filter_banks_9[13] = 32'h00000000;
assign filter_banks_9[14] = 32'h00000000;
assign filter_banks_9[15] = 32'h00000000;
assign filter_banks_9[16] = 32'h00000000;
assign filter_banks_9[17] = 32'h00000000;
assign filter_banks_9[18] = 32'h00000000;
assign filter_banks_9[19] = 32'h00000000;
assign filter_banks_9[20] = 32'h00000000;
assign filter_banks_9[21] = 32'h00000000;
assign filter_banks_9[22] = 32'h00000000;
assign filter_banks_9[23] = 32'h00000000;
assign filter_banks_9[24] = 32'h00000000;
assign filter_banks_9[25] = 32'h3e4ccccd;
assign filter_banks_9[26] = 32'h3ecccccd;
assign filter_banks_9[27] = 32'h3f19999a;
assign filter_banks_9[28] = 32'h3f4ccccd;
assign filter_banks_9[29] = 32'h3f800000;
assign filter_banks_9[30] = 32'h3f4ccccd;
assign filter_banks_9[31] = 32'h3f19999a;
assign filter_banks_9[32] = 32'h3ecccccd;
assign filter_banks_9[33] = 32'h3e4ccccd;
assign filter_banks_9[34] = 32'h00000000;
assign filter_banks_9[35] = 32'h00000000;
assign filter_banks_9[36] = 32'h00000000;
assign filter_banks_9[37] = 32'h00000000;
assign filter_banks_9[38] = 32'h00000000;
assign filter_banks_9[39] = 32'h00000000;
assign filter_banks_9[40] = 32'h00000000;
assign filter_banks_9[41] = 32'h00000000;
assign filter_banks_9[42] = 32'h00000000;
assign filter_banks_9[43] = 32'h00000000;
assign filter_banks_9[44] = 32'h00000000;
assign filter_banks_9[45] = 32'h00000000;
assign filter_banks_9[46] = 32'h00000000;
assign filter_banks_9[47] = 32'h00000000;
assign filter_banks_9[48] = 32'h00000000;
assign filter_banks_9[49] = 32'h00000000;
assign filter_banks_9[50] = 32'h00000000;
assign filter_banks_9[51] = 32'h00000000;
assign filter_banks_9[52] = 32'h00000000;
assign filter_banks_9[53] = 32'h00000000;
assign filter_banks_9[54] = 32'h00000000;
assign filter_banks_9[55] = 32'h00000000;
assign filter_banks_9[56] = 32'h00000000;
assign filter_banks_9[57] = 32'h00000000;
assign filter_banks_9[58] = 32'h00000000;
assign filter_banks_9[59] = 32'h00000000;
assign filter_banks_9[60] = 32'h00000000;
assign filter_banks_9[61] = 32'h00000000;
assign filter_banks_9[62] = 32'h00000000;
assign filter_banks_9[63] = 32'h00000000;
assign filter_banks_9[64] = 32'h00000000;
assign filter_banks_9[65] = 32'h00000000;
assign filter_banks_9[66] = 32'h00000000;
assign filter_banks_9[67] = 32'h00000000;
assign filter_banks_9[68] = 32'h00000000;
assign filter_banks_9[69] = 32'h00000000;
assign filter_banks_9[70] = 32'h00000000;
assign filter_banks_9[71] = 32'h00000000;
assign filter_banks_9[72] = 32'h00000000;
assign filter_banks_9[73] = 32'h00000000;
assign filter_banks_9[74] = 32'h00000000;
assign filter_banks_9[75] = 32'h00000000;
assign filter_banks_9[76] = 32'h00000000;
assign filter_banks_9[77] = 32'h00000000;
assign filter_banks_9[78] = 32'h00000000;
assign filter_banks_9[79] = 32'h00000000;
assign filter_banks_9[80] = 32'h00000000;
assign filter_banks_9[81] = 32'h00000000;
assign filter_banks_9[82] = 32'h00000000;
assign filter_banks_9[83] = 32'h00000000;
assign filter_banks_9[84] = 32'h00000000;
assign filter_banks_9[85] = 32'h00000000;
assign filter_banks_9[86] = 32'h00000000;
assign filter_banks_9[87] = 32'h00000000;
assign filter_banks_9[88] = 32'h00000000;
assign filter_banks_9[89] = 32'h00000000;
assign filter_banks_9[90] = 32'h00000000;
assign filter_banks_9[91] = 32'h00000000;
assign filter_banks_9[92] = 32'h00000000;
assign filter_banks_9[93] = 32'h00000000;
assign filter_banks_9[94] = 32'h00000000;
assign filter_banks_9[95] = 32'h00000000;
assign filter_banks_9[96] = 32'h00000000;
assign filter_banks_9[97] = 32'h00000000;
assign filter_banks_9[98] = 32'h00000000;
assign filter_banks_9[99] = 32'h00000000;
assign filter_banks_9[100] = 32'h00000000;
assign filter_banks_9[101] = 32'h00000000;
assign filter_banks_9[102] = 32'h00000000;
assign filter_banks_9[103] = 32'h00000000;
assign filter_banks_9[104] = 32'h00000000;
assign filter_banks_9[105] = 32'h00000000;
assign filter_banks_9[106] = 32'h00000000;
assign filter_banks_9[107] = 32'h00000000;
assign filter_banks_9[108] = 32'h00000000;
assign filter_banks_9[109] = 32'h00000000;
assign filter_banks_9[110] = 32'h00000000;
assign filter_banks_9[111] = 32'h00000000;
assign filter_banks_9[112] = 32'h00000000;
assign filter_banks_9[113] = 32'h00000000;
assign filter_banks_9[114] = 32'h00000000;
assign filter_banks_9[115] = 32'h00000000;
assign filter_banks_9[116] = 32'h00000000;
assign filter_banks_9[117] = 32'h00000000;
assign filter_banks_9[118] = 32'h00000000;
assign filter_banks_9[119] = 32'h00000000;
assign filter_banks_9[120] = 32'h00000000;
assign filter_banks_9[121] = 32'h00000000;
assign filter_banks_9[122] = 32'h00000000;
assign filter_banks_9[123] = 32'h00000000;
assign filter_banks_9[124] = 32'h00000000;
assign filter_banks_9[125] = 32'h00000000;
assign filter_banks_9[126] = 32'h00000000;
assign filter_banks_9[127] = 32'h00000000;
assign filter_banks_9[128] = 32'h00000000;
assign filter_banks_9[129] = 32'h00000000;
assign filter_banks_9[130] = 32'h00000000;
assign filter_banks_9[131] = 32'h00000000;
assign filter_banks_9[132] = 32'h00000000;
assign filter_banks_9[133] = 32'h00000000;
assign filter_banks_9[134] = 32'h00000000;
assign filter_banks_9[135] = 32'h00000000;
assign filter_banks_9[136] = 32'h00000000;
assign filter_banks_9[137] = 32'h00000000;
assign filter_banks_9[138] = 32'h00000000;
assign filter_banks_9[139] = 32'h00000000;
assign filter_banks_9[140] = 32'h00000000;
assign filter_banks_9[141] = 32'h00000000;
assign filter_banks_9[142] = 32'h00000000;
assign filter_banks_9[143] = 32'h00000000;
assign filter_banks_9[144] = 32'h00000000;
assign filter_banks_9[145] = 32'h00000000;
assign filter_banks_9[146] = 32'h00000000;
assign filter_banks_9[147] = 32'h00000000;
assign filter_banks_9[148] = 32'h00000000;
assign filter_banks_9[149] = 32'h00000000;
assign filter_banks_9[150] = 32'h00000000;
assign filter_banks_9[151] = 32'h00000000;
assign filter_banks_9[152] = 32'h00000000;
assign filter_banks_9[153] = 32'h00000000;
assign filter_banks_9[154] = 32'h00000000;
assign filter_banks_9[155] = 32'h00000000;
assign filter_banks_9[156] = 32'h00000000;
assign filter_banks_9[157] = 32'h00000000;
assign filter_banks_9[158] = 32'h00000000;
assign filter_banks_9[159] = 32'h00000000;
assign filter_banks_9[160] = 32'h00000000;
assign filter_banks_9[161] = 32'h00000000;
assign filter_banks_9[162] = 32'h00000000;
assign filter_banks_9[163] = 32'h00000000;
assign filter_banks_9[164] = 32'h00000000;
assign filter_banks_9[165] = 32'h00000000;
assign filter_banks_9[166] = 32'h00000000;
assign filter_banks_9[167] = 32'h00000000;
assign filter_banks_9[168] = 32'h00000000;
assign filter_banks_9[169] = 32'h00000000;
assign filter_banks_9[170] = 32'h00000000;
assign filter_banks_9[171] = 32'h00000000;
assign filter_banks_9[172] = 32'h00000000;
assign filter_banks_9[173] = 32'h00000000;
assign filter_banks_9[174] = 32'h00000000;
assign filter_banks_9[175] = 32'h00000000;
assign filter_banks_9[176] = 32'h00000000;
assign filter_banks_9[177] = 32'h00000000;
assign filter_banks_9[178] = 32'h00000000;
assign filter_banks_9[179] = 32'h00000000;
assign filter_banks_9[180] = 32'h00000000;
assign filter_banks_9[181] = 32'h00000000;
assign filter_banks_9[182] = 32'h00000000;
assign filter_banks_9[183] = 32'h00000000;
assign filter_banks_9[184] = 32'h00000000;
assign filter_banks_9[185] = 32'h00000000;
assign filter_banks_9[186] = 32'h00000000;
assign filter_banks_9[187] = 32'h00000000;
assign filter_banks_9[188] = 32'h00000000;
assign filter_banks_9[189] = 32'h00000000;
assign filter_banks_9[190] = 32'h00000000;
assign filter_banks_9[191] = 32'h00000000;
assign filter_banks_9[192] = 32'h00000000;
assign filter_banks_9[193] = 32'h00000000;
assign filter_banks_9[194] = 32'h00000000;
assign filter_banks_9[195] = 32'h00000000;
assign filter_banks_9[196] = 32'h00000000;
assign filter_banks_9[197] = 32'h00000000;
assign filter_banks_9[198] = 32'h00000000;
assign filter_banks_9[199] = 32'h00000000;
assign filter_banks_9[200] = 32'h00000000;
assign filter_banks_9[201] = 32'h00000000;
assign filter_banks_9[202] = 32'h00000000;
assign filter_banks_9[203] = 32'h00000000;
assign filter_banks_9[204] = 32'h00000000;
assign filter_banks_9[205] = 32'h00000000;
assign filter_banks_9[206] = 32'h00000000;
assign filter_banks_9[207] = 32'h00000000;
assign filter_banks_9[208] = 32'h00000000;
assign filter_banks_9[209] = 32'h00000000;
assign filter_banks_9[210] = 32'h00000000;
assign filter_banks_9[211] = 32'h00000000;
assign filter_banks_9[212] = 32'h00000000;
assign filter_banks_9[213] = 32'h00000000;
assign filter_banks_9[214] = 32'h00000000;
assign filter_banks_9[215] = 32'h00000000;
assign filter_banks_9[216] = 32'h00000000;
assign filter_banks_9[217] = 32'h00000000;
assign filter_banks_9[218] = 32'h00000000;
assign filter_banks_9[219] = 32'h00000000;
assign filter_banks_9[220] = 32'h00000000;
assign filter_banks_9[221] = 32'h00000000;
assign filter_banks_9[222] = 32'h00000000;
assign filter_banks_9[223] = 32'h00000000;
assign filter_banks_9[224] = 32'h00000000;
assign filter_banks_9[225] = 32'h00000000;
assign filter_banks_9[226] = 32'h00000000;
assign filter_banks_9[227] = 32'h00000000;
assign filter_banks_9[228] = 32'h00000000;
assign filter_banks_9[229] = 32'h00000000;
assign filter_banks_9[230] = 32'h00000000;
assign filter_banks_9[231] = 32'h00000000;
assign filter_banks_9[232] = 32'h00000000;
assign filter_banks_9[233] = 32'h00000000;
assign filter_banks_9[234] = 32'h00000000;
assign filter_banks_9[235] = 32'h00000000;
assign filter_banks_9[236] = 32'h00000000;
assign filter_banks_9[237] = 32'h00000000;
assign filter_banks_9[238] = 32'h00000000;
assign filter_banks_9[239] = 32'h00000000;
assign filter_banks_9[240] = 32'h00000000;
assign filter_banks_9[241] = 32'h00000000;
assign filter_banks_9[242] = 32'h00000000;
assign filter_banks_9[243] = 32'h00000000;
assign filter_banks_9[244] = 32'h00000000;
assign filter_banks_9[245] = 32'h00000000;
assign filter_banks_9[246] = 32'h00000000;
assign filter_banks_9[247] = 32'h00000000;
assign filter_banks_9[248] = 32'h00000000;
assign filter_banks_9[249] = 32'h00000000;
assign filter_banks_9[250] = 32'h00000000;
assign filter_banks_9[251] = 32'h00000000;
assign filter_banks_9[252] = 32'h00000000;
assign filter_banks_9[253] = 32'h00000000;
assign filter_banks_9[254] = 32'h00000000;
assign filter_banks_9[255] = 32'h00000000;
assign filter_banks_9[256] = 32'h00000000;
assign filter_banks_10[0] = 32'h00000000;
assign filter_banks_10[1] = 32'h00000000;
assign filter_banks_10[2] = 32'h00000000;
assign filter_banks_10[3] = 32'h00000000;
assign filter_banks_10[4] = 32'h00000000;
assign filter_banks_10[5] = 32'h00000000;
assign filter_banks_10[6] = 32'h00000000;
assign filter_banks_10[7] = 32'h00000000;
assign filter_banks_10[8] = 32'h00000000;
assign filter_banks_10[9] = 32'h00000000;
assign filter_banks_10[10] = 32'h00000000;
assign filter_banks_10[11] = 32'h00000000;
assign filter_banks_10[12] = 32'h00000000;
assign filter_banks_10[13] = 32'h00000000;
assign filter_banks_10[14] = 32'h00000000;
assign filter_banks_10[15] = 32'h00000000;
assign filter_banks_10[16] = 32'h00000000;
assign filter_banks_10[17] = 32'h00000000;
assign filter_banks_10[18] = 32'h00000000;
assign filter_banks_10[19] = 32'h00000000;
assign filter_banks_10[20] = 32'h00000000;
assign filter_banks_10[21] = 32'h00000000;
assign filter_banks_10[22] = 32'h00000000;
assign filter_banks_10[23] = 32'h00000000;
assign filter_banks_10[24] = 32'h00000000;
assign filter_banks_10[25] = 32'h00000000;
assign filter_banks_10[26] = 32'h00000000;
assign filter_banks_10[27] = 32'h00000000;
assign filter_banks_10[28] = 32'h00000000;
assign filter_banks_10[29] = 32'h00000000;
assign filter_banks_10[30] = 32'h3e4ccccd;
assign filter_banks_10[31] = 32'h3ecccccd;
assign filter_banks_10[32] = 32'h3f19999a;
assign filter_banks_10[33] = 32'h3f4ccccd;
assign filter_banks_10[34] = 32'h3f800000;
assign filter_banks_10[35] = 32'h3f555555;
assign filter_banks_10[36] = 32'h3f2aaaab;
assign filter_banks_10[37] = 32'h3f000000;
assign filter_banks_10[38] = 32'h3eaaaaab;
assign filter_banks_10[39] = 32'h3e2aaaab;
assign filter_banks_10[40] = 32'h00000000;
assign filter_banks_10[41] = 32'h00000000;
assign filter_banks_10[42] = 32'h00000000;
assign filter_banks_10[43] = 32'h00000000;
assign filter_banks_10[44] = 32'h00000000;
assign filter_banks_10[45] = 32'h00000000;
assign filter_banks_10[46] = 32'h00000000;
assign filter_banks_10[47] = 32'h00000000;
assign filter_banks_10[48] = 32'h00000000;
assign filter_banks_10[49] = 32'h00000000;
assign filter_banks_10[50] = 32'h00000000;
assign filter_banks_10[51] = 32'h00000000;
assign filter_banks_10[52] = 32'h00000000;
assign filter_banks_10[53] = 32'h00000000;
assign filter_banks_10[54] = 32'h00000000;
assign filter_banks_10[55] = 32'h00000000;
assign filter_banks_10[56] = 32'h00000000;
assign filter_banks_10[57] = 32'h00000000;
assign filter_banks_10[58] = 32'h00000000;
assign filter_banks_10[59] = 32'h00000000;
assign filter_banks_10[60] = 32'h00000000;
assign filter_banks_10[61] = 32'h00000000;
assign filter_banks_10[62] = 32'h00000000;
assign filter_banks_10[63] = 32'h00000000;
assign filter_banks_10[64] = 32'h00000000;
assign filter_banks_10[65] = 32'h00000000;
assign filter_banks_10[66] = 32'h00000000;
assign filter_banks_10[67] = 32'h00000000;
assign filter_banks_10[68] = 32'h00000000;
assign filter_banks_10[69] = 32'h00000000;
assign filter_banks_10[70] = 32'h00000000;
assign filter_banks_10[71] = 32'h00000000;
assign filter_banks_10[72] = 32'h00000000;
assign filter_banks_10[73] = 32'h00000000;
assign filter_banks_10[74] = 32'h00000000;
assign filter_banks_10[75] = 32'h00000000;
assign filter_banks_10[76] = 32'h00000000;
assign filter_banks_10[77] = 32'h00000000;
assign filter_banks_10[78] = 32'h00000000;
assign filter_banks_10[79] = 32'h00000000;
assign filter_banks_10[80] = 32'h00000000;
assign filter_banks_10[81] = 32'h00000000;
assign filter_banks_10[82] = 32'h00000000;
assign filter_banks_10[83] = 32'h00000000;
assign filter_banks_10[84] = 32'h00000000;
assign filter_banks_10[85] = 32'h00000000;
assign filter_banks_10[86] = 32'h00000000;
assign filter_banks_10[87] = 32'h00000000;
assign filter_banks_10[88] = 32'h00000000;
assign filter_banks_10[89] = 32'h00000000;
assign filter_banks_10[90] = 32'h00000000;
assign filter_banks_10[91] = 32'h00000000;
assign filter_banks_10[92] = 32'h00000000;
assign filter_banks_10[93] = 32'h00000000;
assign filter_banks_10[94] = 32'h00000000;
assign filter_banks_10[95] = 32'h00000000;
assign filter_banks_10[96] = 32'h00000000;
assign filter_banks_10[97] = 32'h00000000;
assign filter_banks_10[98] = 32'h00000000;
assign filter_banks_10[99] = 32'h00000000;
assign filter_banks_10[100] = 32'h00000000;
assign filter_banks_10[101] = 32'h00000000;
assign filter_banks_10[102] = 32'h00000000;
assign filter_banks_10[103] = 32'h00000000;
assign filter_banks_10[104] = 32'h00000000;
assign filter_banks_10[105] = 32'h00000000;
assign filter_banks_10[106] = 32'h00000000;
assign filter_banks_10[107] = 32'h00000000;
assign filter_banks_10[108] = 32'h00000000;
assign filter_banks_10[109] = 32'h00000000;
assign filter_banks_10[110] = 32'h00000000;
assign filter_banks_10[111] = 32'h00000000;
assign filter_banks_10[112] = 32'h00000000;
assign filter_banks_10[113] = 32'h00000000;
assign filter_banks_10[114] = 32'h00000000;
assign filter_banks_10[115] = 32'h00000000;
assign filter_banks_10[116] = 32'h00000000;
assign filter_banks_10[117] = 32'h00000000;
assign filter_banks_10[118] = 32'h00000000;
assign filter_banks_10[119] = 32'h00000000;
assign filter_banks_10[120] = 32'h00000000;
assign filter_banks_10[121] = 32'h00000000;
assign filter_banks_10[122] = 32'h00000000;
assign filter_banks_10[123] = 32'h00000000;
assign filter_banks_10[124] = 32'h00000000;
assign filter_banks_10[125] = 32'h00000000;
assign filter_banks_10[126] = 32'h00000000;
assign filter_banks_10[127] = 32'h00000000;
assign filter_banks_10[128] = 32'h00000000;
assign filter_banks_10[129] = 32'h00000000;
assign filter_banks_10[130] = 32'h00000000;
assign filter_banks_10[131] = 32'h00000000;
assign filter_banks_10[132] = 32'h00000000;
assign filter_banks_10[133] = 32'h00000000;
assign filter_banks_10[134] = 32'h00000000;
assign filter_banks_10[135] = 32'h00000000;
assign filter_banks_10[136] = 32'h00000000;
assign filter_banks_10[137] = 32'h00000000;
assign filter_banks_10[138] = 32'h00000000;
assign filter_banks_10[139] = 32'h00000000;
assign filter_banks_10[140] = 32'h00000000;
assign filter_banks_10[141] = 32'h00000000;
assign filter_banks_10[142] = 32'h00000000;
assign filter_banks_10[143] = 32'h00000000;
assign filter_banks_10[144] = 32'h00000000;
assign filter_banks_10[145] = 32'h00000000;
assign filter_banks_10[146] = 32'h00000000;
assign filter_banks_10[147] = 32'h00000000;
assign filter_banks_10[148] = 32'h00000000;
assign filter_banks_10[149] = 32'h00000000;
assign filter_banks_10[150] = 32'h00000000;
assign filter_banks_10[151] = 32'h00000000;
assign filter_banks_10[152] = 32'h00000000;
assign filter_banks_10[153] = 32'h00000000;
assign filter_banks_10[154] = 32'h00000000;
assign filter_banks_10[155] = 32'h00000000;
assign filter_banks_10[156] = 32'h00000000;
assign filter_banks_10[157] = 32'h00000000;
assign filter_banks_10[158] = 32'h00000000;
assign filter_banks_10[159] = 32'h00000000;
assign filter_banks_10[160] = 32'h00000000;
assign filter_banks_10[161] = 32'h00000000;
assign filter_banks_10[162] = 32'h00000000;
assign filter_banks_10[163] = 32'h00000000;
assign filter_banks_10[164] = 32'h00000000;
assign filter_banks_10[165] = 32'h00000000;
assign filter_banks_10[166] = 32'h00000000;
assign filter_banks_10[167] = 32'h00000000;
assign filter_banks_10[168] = 32'h00000000;
assign filter_banks_10[169] = 32'h00000000;
assign filter_banks_10[170] = 32'h00000000;
assign filter_banks_10[171] = 32'h00000000;
assign filter_banks_10[172] = 32'h00000000;
assign filter_banks_10[173] = 32'h00000000;
assign filter_banks_10[174] = 32'h00000000;
assign filter_banks_10[175] = 32'h00000000;
assign filter_banks_10[176] = 32'h00000000;
assign filter_banks_10[177] = 32'h00000000;
assign filter_banks_10[178] = 32'h00000000;
assign filter_banks_10[179] = 32'h00000000;
assign filter_banks_10[180] = 32'h00000000;
assign filter_banks_10[181] = 32'h00000000;
assign filter_banks_10[182] = 32'h00000000;
assign filter_banks_10[183] = 32'h00000000;
assign filter_banks_10[184] = 32'h00000000;
assign filter_banks_10[185] = 32'h00000000;
assign filter_banks_10[186] = 32'h00000000;
assign filter_banks_10[187] = 32'h00000000;
assign filter_banks_10[188] = 32'h00000000;
assign filter_banks_10[189] = 32'h00000000;
assign filter_banks_10[190] = 32'h00000000;
assign filter_banks_10[191] = 32'h00000000;
assign filter_banks_10[192] = 32'h00000000;
assign filter_banks_10[193] = 32'h00000000;
assign filter_banks_10[194] = 32'h00000000;
assign filter_banks_10[195] = 32'h00000000;
assign filter_banks_10[196] = 32'h00000000;
assign filter_banks_10[197] = 32'h00000000;
assign filter_banks_10[198] = 32'h00000000;
assign filter_banks_10[199] = 32'h00000000;
assign filter_banks_10[200] = 32'h00000000;
assign filter_banks_10[201] = 32'h00000000;
assign filter_banks_10[202] = 32'h00000000;
assign filter_banks_10[203] = 32'h00000000;
assign filter_banks_10[204] = 32'h00000000;
assign filter_banks_10[205] = 32'h00000000;
assign filter_banks_10[206] = 32'h00000000;
assign filter_banks_10[207] = 32'h00000000;
assign filter_banks_10[208] = 32'h00000000;
assign filter_banks_10[209] = 32'h00000000;
assign filter_banks_10[210] = 32'h00000000;
assign filter_banks_10[211] = 32'h00000000;
assign filter_banks_10[212] = 32'h00000000;
assign filter_banks_10[213] = 32'h00000000;
assign filter_banks_10[214] = 32'h00000000;
assign filter_banks_10[215] = 32'h00000000;
assign filter_banks_10[216] = 32'h00000000;
assign filter_banks_10[217] = 32'h00000000;
assign filter_banks_10[218] = 32'h00000000;
assign filter_banks_10[219] = 32'h00000000;
assign filter_banks_10[220] = 32'h00000000;
assign filter_banks_10[221] = 32'h00000000;
assign filter_banks_10[222] = 32'h00000000;
assign filter_banks_10[223] = 32'h00000000;
assign filter_banks_10[224] = 32'h00000000;
assign filter_banks_10[225] = 32'h00000000;
assign filter_banks_10[226] = 32'h00000000;
assign filter_banks_10[227] = 32'h00000000;
assign filter_banks_10[228] = 32'h00000000;
assign filter_banks_10[229] = 32'h00000000;
assign filter_banks_10[230] = 32'h00000000;
assign filter_banks_10[231] = 32'h00000000;
assign filter_banks_10[232] = 32'h00000000;
assign filter_banks_10[233] = 32'h00000000;
assign filter_banks_10[234] = 32'h00000000;
assign filter_banks_10[235] = 32'h00000000;
assign filter_banks_10[236] = 32'h00000000;
assign filter_banks_10[237] = 32'h00000000;
assign filter_banks_10[238] = 32'h00000000;
assign filter_banks_10[239] = 32'h00000000;
assign filter_banks_10[240] = 32'h00000000;
assign filter_banks_10[241] = 32'h00000000;
assign filter_banks_10[242] = 32'h00000000;
assign filter_banks_10[243] = 32'h00000000;
assign filter_banks_10[244] = 32'h00000000;
assign filter_banks_10[245] = 32'h00000000;
assign filter_banks_10[246] = 32'h00000000;
assign filter_banks_10[247] = 32'h00000000;
assign filter_banks_10[248] = 32'h00000000;
assign filter_banks_10[249] = 32'h00000000;
assign filter_banks_10[250] = 32'h00000000;
assign filter_banks_10[251] = 32'h00000000;
assign filter_banks_10[252] = 32'h00000000;
assign filter_banks_10[253] = 32'h00000000;
assign filter_banks_10[254] = 32'h00000000;
assign filter_banks_10[255] = 32'h00000000;
assign filter_banks_10[256] = 32'h00000000;
assign filter_banks_11[0] = 32'h00000000;
assign filter_banks_11[1] = 32'h00000000;
assign filter_banks_11[2] = 32'h00000000;
assign filter_banks_11[3] = 32'h00000000;
assign filter_banks_11[4] = 32'h00000000;
assign filter_banks_11[5] = 32'h00000000;
assign filter_banks_11[6] = 32'h00000000;
assign filter_banks_11[7] = 32'h00000000;
assign filter_banks_11[8] = 32'h00000000;
assign filter_banks_11[9] = 32'h00000000;
assign filter_banks_11[10] = 32'h00000000;
assign filter_banks_11[11] = 32'h00000000;
assign filter_banks_11[12] = 32'h00000000;
assign filter_banks_11[13] = 32'h00000000;
assign filter_banks_11[14] = 32'h00000000;
assign filter_banks_11[15] = 32'h00000000;
assign filter_banks_11[16] = 32'h00000000;
assign filter_banks_11[17] = 32'h00000000;
assign filter_banks_11[18] = 32'h00000000;
assign filter_banks_11[19] = 32'h00000000;
assign filter_banks_11[20] = 32'h00000000;
assign filter_banks_11[21] = 32'h00000000;
assign filter_banks_11[22] = 32'h00000000;
assign filter_banks_11[23] = 32'h00000000;
assign filter_banks_11[24] = 32'h00000000;
assign filter_banks_11[25] = 32'h00000000;
assign filter_banks_11[26] = 32'h00000000;
assign filter_banks_11[27] = 32'h00000000;
assign filter_banks_11[28] = 32'h00000000;
assign filter_banks_11[29] = 32'h00000000;
assign filter_banks_11[30] = 32'h00000000;
assign filter_banks_11[31] = 32'h00000000;
assign filter_banks_11[32] = 32'h00000000;
assign filter_banks_11[33] = 32'h00000000;
assign filter_banks_11[34] = 32'h00000000;
assign filter_banks_11[35] = 32'h3e2aaaab;
assign filter_banks_11[36] = 32'h3eaaaaab;
assign filter_banks_11[37] = 32'h3f000000;
assign filter_banks_11[38] = 32'h3f2aaaab;
assign filter_banks_11[39] = 32'h3f555555;
assign filter_banks_11[40] = 32'h3f800000;
assign filter_banks_11[41] = 32'h3f555555;
assign filter_banks_11[42] = 32'h3f2aaaab;
assign filter_banks_11[43] = 32'h3f000000;
assign filter_banks_11[44] = 32'h3eaaaaab;
assign filter_banks_11[45] = 32'h3e2aaaab;
assign filter_banks_11[46] = 32'h00000000;
assign filter_banks_11[47] = 32'h00000000;
assign filter_banks_11[48] = 32'h00000000;
assign filter_banks_11[49] = 32'h00000000;
assign filter_banks_11[50] = 32'h00000000;
assign filter_banks_11[51] = 32'h00000000;
assign filter_banks_11[52] = 32'h00000000;
assign filter_banks_11[53] = 32'h00000000;
assign filter_banks_11[54] = 32'h00000000;
assign filter_banks_11[55] = 32'h00000000;
assign filter_banks_11[56] = 32'h00000000;
assign filter_banks_11[57] = 32'h00000000;
assign filter_banks_11[58] = 32'h00000000;
assign filter_banks_11[59] = 32'h00000000;
assign filter_banks_11[60] = 32'h00000000;
assign filter_banks_11[61] = 32'h00000000;
assign filter_banks_11[62] = 32'h00000000;
assign filter_banks_11[63] = 32'h00000000;
assign filter_banks_11[64] = 32'h00000000;
assign filter_banks_11[65] = 32'h00000000;
assign filter_banks_11[66] = 32'h00000000;
assign filter_banks_11[67] = 32'h00000000;
assign filter_banks_11[68] = 32'h00000000;
assign filter_banks_11[69] = 32'h00000000;
assign filter_banks_11[70] = 32'h00000000;
assign filter_banks_11[71] = 32'h00000000;
assign filter_banks_11[72] = 32'h00000000;
assign filter_banks_11[73] = 32'h00000000;
assign filter_banks_11[74] = 32'h00000000;
assign filter_banks_11[75] = 32'h00000000;
assign filter_banks_11[76] = 32'h00000000;
assign filter_banks_11[77] = 32'h00000000;
assign filter_banks_11[78] = 32'h00000000;
assign filter_banks_11[79] = 32'h00000000;
assign filter_banks_11[80] = 32'h00000000;
assign filter_banks_11[81] = 32'h00000000;
assign filter_banks_11[82] = 32'h00000000;
assign filter_banks_11[83] = 32'h00000000;
assign filter_banks_11[84] = 32'h00000000;
assign filter_banks_11[85] = 32'h00000000;
assign filter_banks_11[86] = 32'h00000000;
assign filter_banks_11[87] = 32'h00000000;
assign filter_banks_11[88] = 32'h00000000;
assign filter_banks_11[89] = 32'h00000000;
assign filter_banks_11[90] = 32'h00000000;
assign filter_banks_11[91] = 32'h00000000;
assign filter_banks_11[92] = 32'h00000000;
assign filter_banks_11[93] = 32'h00000000;
assign filter_banks_11[94] = 32'h00000000;
assign filter_banks_11[95] = 32'h00000000;
assign filter_banks_11[96] = 32'h00000000;
assign filter_banks_11[97] = 32'h00000000;
assign filter_banks_11[98] = 32'h00000000;
assign filter_banks_11[99] = 32'h00000000;
assign filter_banks_11[100] = 32'h00000000;
assign filter_banks_11[101] = 32'h00000000;
assign filter_banks_11[102] = 32'h00000000;
assign filter_banks_11[103] = 32'h00000000;
assign filter_banks_11[104] = 32'h00000000;
assign filter_banks_11[105] = 32'h00000000;
assign filter_banks_11[106] = 32'h00000000;
assign filter_banks_11[107] = 32'h00000000;
assign filter_banks_11[108] = 32'h00000000;
assign filter_banks_11[109] = 32'h00000000;
assign filter_banks_11[110] = 32'h00000000;
assign filter_banks_11[111] = 32'h00000000;
assign filter_banks_11[112] = 32'h00000000;
assign filter_banks_11[113] = 32'h00000000;
assign filter_banks_11[114] = 32'h00000000;
assign filter_banks_11[115] = 32'h00000000;
assign filter_banks_11[116] = 32'h00000000;
assign filter_banks_11[117] = 32'h00000000;
assign filter_banks_11[118] = 32'h00000000;
assign filter_banks_11[119] = 32'h00000000;
assign filter_banks_11[120] = 32'h00000000;
assign filter_banks_11[121] = 32'h00000000;
assign filter_banks_11[122] = 32'h00000000;
assign filter_banks_11[123] = 32'h00000000;
assign filter_banks_11[124] = 32'h00000000;
assign filter_banks_11[125] = 32'h00000000;
assign filter_banks_11[126] = 32'h00000000;
assign filter_banks_11[127] = 32'h00000000;
assign filter_banks_11[128] = 32'h00000000;
assign filter_banks_11[129] = 32'h00000000;
assign filter_banks_11[130] = 32'h00000000;
assign filter_banks_11[131] = 32'h00000000;
assign filter_banks_11[132] = 32'h00000000;
assign filter_banks_11[133] = 32'h00000000;
assign filter_banks_11[134] = 32'h00000000;
assign filter_banks_11[135] = 32'h00000000;
assign filter_banks_11[136] = 32'h00000000;
assign filter_banks_11[137] = 32'h00000000;
assign filter_banks_11[138] = 32'h00000000;
assign filter_banks_11[139] = 32'h00000000;
assign filter_banks_11[140] = 32'h00000000;
assign filter_banks_11[141] = 32'h00000000;
assign filter_banks_11[142] = 32'h00000000;
assign filter_banks_11[143] = 32'h00000000;
assign filter_banks_11[144] = 32'h00000000;
assign filter_banks_11[145] = 32'h00000000;
assign filter_banks_11[146] = 32'h00000000;
assign filter_banks_11[147] = 32'h00000000;
assign filter_banks_11[148] = 32'h00000000;
assign filter_banks_11[149] = 32'h00000000;
assign filter_banks_11[150] = 32'h00000000;
assign filter_banks_11[151] = 32'h00000000;
assign filter_banks_11[152] = 32'h00000000;
assign filter_banks_11[153] = 32'h00000000;
assign filter_banks_11[154] = 32'h00000000;
assign filter_banks_11[155] = 32'h00000000;
assign filter_banks_11[156] = 32'h00000000;
assign filter_banks_11[157] = 32'h00000000;
assign filter_banks_11[158] = 32'h00000000;
assign filter_banks_11[159] = 32'h00000000;
assign filter_banks_11[160] = 32'h00000000;
assign filter_banks_11[161] = 32'h00000000;
assign filter_banks_11[162] = 32'h00000000;
assign filter_banks_11[163] = 32'h00000000;
assign filter_banks_11[164] = 32'h00000000;
assign filter_banks_11[165] = 32'h00000000;
assign filter_banks_11[166] = 32'h00000000;
assign filter_banks_11[167] = 32'h00000000;
assign filter_banks_11[168] = 32'h00000000;
assign filter_banks_11[169] = 32'h00000000;
assign filter_banks_11[170] = 32'h00000000;
assign filter_banks_11[171] = 32'h00000000;
assign filter_banks_11[172] = 32'h00000000;
assign filter_banks_11[173] = 32'h00000000;
assign filter_banks_11[174] = 32'h00000000;
assign filter_banks_11[175] = 32'h00000000;
assign filter_banks_11[176] = 32'h00000000;
assign filter_banks_11[177] = 32'h00000000;
assign filter_banks_11[178] = 32'h00000000;
assign filter_banks_11[179] = 32'h00000000;
assign filter_banks_11[180] = 32'h00000000;
assign filter_banks_11[181] = 32'h00000000;
assign filter_banks_11[182] = 32'h00000000;
assign filter_banks_11[183] = 32'h00000000;
assign filter_banks_11[184] = 32'h00000000;
assign filter_banks_11[185] = 32'h00000000;
assign filter_banks_11[186] = 32'h00000000;
assign filter_banks_11[187] = 32'h00000000;
assign filter_banks_11[188] = 32'h00000000;
assign filter_banks_11[189] = 32'h00000000;
assign filter_banks_11[190] = 32'h00000000;
assign filter_banks_11[191] = 32'h00000000;
assign filter_banks_11[192] = 32'h00000000;
assign filter_banks_11[193] = 32'h00000000;
assign filter_banks_11[194] = 32'h00000000;
assign filter_banks_11[195] = 32'h00000000;
assign filter_banks_11[196] = 32'h00000000;
assign filter_banks_11[197] = 32'h00000000;
assign filter_banks_11[198] = 32'h00000000;
assign filter_banks_11[199] = 32'h00000000;
assign filter_banks_11[200] = 32'h00000000;
assign filter_banks_11[201] = 32'h00000000;
assign filter_banks_11[202] = 32'h00000000;
assign filter_banks_11[203] = 32'h00000000;
assign filter_banks_11[204] = 32'h00000000;
assign filter_banks_11[205] = 32'h00000000;
assign filter_banks_11[206] = 32'h00000000;
assign filter_banks_11[207] = 32'h00000000;
assign filter_banks_11[208] = 32'h00000000;
assign filter_banks_11[209] = 32'h00000000;
assign filter_banks_11[210] = 32'h00000000;
assign filter_banks_11[211] = 32'h00000000;
assign filter_banks_11[212] = 32'h00000000;
assign filter_banks_11[213] = 32'h00000000;
assign filter_banks_11[214] = 32'h00000000;
assign filter_banks_11[215] = 32'h00000000;
assign filter_banks_11[216] = 32'h00000000;
assign filter_banks_11[217] = 32'h00000000;
assign filter_banks_11[218] = 32'h00000000;
assign filter_banks_11[219] = 32'h00000000;
assign filter_banks_11[220] = 32'h00000000;
assign filter_banks_11[221] = 32'h00000000;
assign filter_banks_11[222] = 32'h00000000;
assign filter_banks_11[223] = 32'h00000000;
assign filter_banks_11[224] = 32'h00000000;
assign filter_banks_11[225] = 32'h00000000;
assign filter_banks_11[226] = 32'h00000000;
assign filter_banks_11[227] = 32'h00000000;
assign filter_banks_11[228] = 32'h00000000;
assign filter_banks_11[229] = 32'h00000000;
assign filter_banks_11[230] = 32'h00000000;
assign filter_banks_11[231] = 32'h00000000;
assign filter_banks_11[232] = 32'h00000000;
assign filter_banks_11[233] = 32'h00000000;
assign filter_banks_11[234] = 32'h00000000;
assign filter_banks_11[235] = 32'h00000000;
assign filter_banks_11[236] = 32'h00000000;
assign filter_banks_11[237] = 32'h00000000;
assign filter_banks_11[238] = 32'h00000000;
assign filter_banks_11[239] = 32'h00000000;
assign filter_banks_11[240] = 32'h00000000;
assign filter_banks_11[241] = 32'h00000000;
assign filter_banks_11[242] = 32'h00000000;
assign filter_banks_11[243] = 32'h00000000;
assign filter_banks_11[244] = 32'h00000000;
assign filter_banks_11[245] = 32'h00000000;
assign filter_banks_11[246] = 32'h00000000;
assign filter_banks_11[247] = 32'h00000000;
assign filter_banks_11[248] = 32'h00000000;
assign filter_banks_11[249] = 32'h00000000;
assign filter_banks_11[250] = 32'h00000000;
assign filter_banks_11[251] = 32'h00000000;
assign filter_banks_11[252] = 32'h00000000;
assign filter_banks_11[253] = 32'h00000000;
assign filter_banks_11[254] = 32'h00000000;
assign filter_banks_11[255] = 32'h00000000;
assign filter_banks_11[256] = 32'h00000000;
assign filter_banks_12[0] = 32'h00000000;
assign filter_banks_12[1] = 32'h00000000;
assign filter_banks_12[2] = 32'h00000000;
assign filter_banks_12[3] = 32'h00000000;
assign filter_banks_12[4] = 32'h00000000;
assign filter_banks_12[5] = 32'h00000000;
assign filter_banks_12[6] = 32'h00000000;
assign filter_banks_12[7] = 32'h00000000;
assign filter_banks_12[8] = 32'h00000000;
assign filter_banks_12[9] = 32'h00000000;
assign filter_banks_12[10] = 32'h00000000;
assign filter_banks_12[11] = 32'h00000000;
assign filter_banks_12[12] = 32'h00000000;
assign filter_banks_12[13] = 32'h00000000;
assign filter_banks_12[14] = 32'h00000000;
assign filter_banks_12[15] = 32'h00000000;
assign filter_banks_12[16] = 32'h00000000;
assign filter_banks_12[17] = 32'h00000000;
assign filter_banks_12[18] = 32'h00000000;
assign filter_banks_12[19] = 32'h00000000;
assign filter_banks_12[20] = 32'h00000000;
assign filter_banks_12[21] = 32'h00000000;
assign filter_banks_12[22] = 32'h00000000;
assign filter_banks_12[23] = 32'h00000000;
assign filter_banks_12[24] = 32'h00000000;
assign filter_banks_12[25] = 32'h00000000;
assign filter_banks_12[26] = 32'h00000000;
assign filter_banks_12[27] = 32'h00000000;
assign filter_banks_12[28] = 32'h00000000;
assign filter_banks_12[29] = 32'h00000000;
assign filter_banks_12[30] = 32'h00000000;
assign filter_banks_12[31] = 32'h00000000;
assign filter_banks_12[32] = 32'h00000000;
assign filter_banks_12[33] = 32'h00000000;
assign filter_banks_12[34] = 32'h00000000;
assign filter_banks_12[35] = 32'h00000000;
assign filter_banks_12[36] = 32'h00000000;
assign filter_banks_12[37] = 32'h00000000;
assign filter_banks_12[38] = 32'h00000000;
assign filter_banks_12[39] = 32'h00000000;
assign filter_banks_12[40] = 32'h00000000;
assign filter_banks_12[41] = 32'h3e2aaaab;
assign filter_banks_12[42] = 32'h3eaaaaab;
assign filter_banks_12[43] = 32'h3f000000;
assign filter_banks_12[44] = 32'h3f2aaaab;
assign filter_banks_12[45] = 32'h3f555555;
assign filter_banks_12[46] = 32'h3f800000;
assign filter_banks_12[47] = 32'h3f5b6db7;
assign filter_banks_12[48] = 32'h3f36db6e;
assign filter_banks_12[49] = 32'h3f124925;
assign filter_banks_12[50] = 32'h3edb6db7;
assign filter_banks_12[51] = 32'h3e924925;
assign filter_banks_12[52] = 32'h3e124925;
assign filter_banks_12[53] = 32'h00000000;
assign filter_banks_12[54] = 32'h00000000;
assign filter_banks_12[55] = 32'h00000000;
assign filter_banks_12[56] = 32'h00000000;
assign filter_banks_12[57] = 32'h00000000;
assign filter_banks_12[58] = 32'h00000000;
assign filter_banks_12[59] = 32'h00000000;
assign filter_banks_12[60] = 32'h00000000;
assign filter_banks_12[61] = 32'h00000000;
assign filter_banks_12[62] = 32'h00000000;
assign filter_banks_12[63] = 32'h00000000;
assign filter_banks_12[64] = 32'h00000000;
assign filter_banks_12[65] = 32'h00000000;
assign filter_banks_12[66] = 32'h00000000;
assign filter_banks_12[67] = 32'h00000000;
assign filter_banks_12[68] = 32'h00000000;
assign filter_banks_12[69] = 32'h00000000;
assign filter_banks_12[70] = 32'h00000000;
assign filter_banks_12[71] = 32'h00000000;
assign filter_banks_12[72] = 32'h00000000;
assign filter_banks_12[73] = 32'h00000000;
assign filter_banks_12[74] = 32'h00000000;
assign filter_banks_12[75] = 32'h00000000;
assign filter_banks_12[76] = 32'h00000000;
assign filter_banks_12[77] = 32'h00000000;
assign filter_banks_12[78] = 32'h00000000;
assign filter_banks_12[79] = 32'h00000000;
assign filter_banks_12[80] = 32'h00000000;
assign filter_banks_12[81] = 32'h00000000;
assign filter_banks_12[82] = 32'h00000000;
assign filter_banks_12[83] = 32'h00000000;
assign filter_banks_12[84] = 32'h00000000;
assign filter_banks_12[85] = 32'h00000000;
assign filter_banks_12[86] = 32'h00000000;
assign filter_banks_12[87] = 32'h00000000;
assign filter_banks_12[88] = 32'h00000000;
assign filter_banks_12[89] = 32'h00000000;
assign filter_banks_12[90] = 32'h00000000;
assign filter_banks_12[91] = 32'h00000000;
assign filter_banks_12[92] = 32'h00000000;
assign filter_banks_12[93] = 32'h00000000;
assign filter_banks_12[94] = 32'h00000000;
assign filter_banks_12[95] = 32'h00000000;
assign filter_banks_12[96] = 32'h00000000;
assign filter_banks_12[97] = 32'h00000000;
assign filter_banks_12[98] = 32'h00000000;
assign filter_banks_12[99] = 32'h00000000;
assign filter_banks_12[100] = 32'h00000000;
assign filter_banks_12[101] = 32'h00000000;
assign filter_banks_12[102] = 32'h00000000;
assign filter_banks_12[103] = 32'h00000000;
assign filter_banks_12[104] = 32'h00000000;
assign filter_banks_12[105] = 32'h00000000;
assign filter_banks_12[106] = 32'h00000000;
assign filter_banks_12[107] = 32'h00000000;
assign filter_banks_12[108] = 32'h00000000;
assign filter_banks_12[109] = 32'h00000000;
assign filter_banks_12[110] = 32'h00000000;
assign filter_banks_12[111] = 32'h00000000;
assign filter_banks_12[112] = 32'h00000000;
assign filter_banks_12[113] = 32'h00000000;
assign filter_banks_12[114] = 32'h00000000;
assign filter_banks_12[115] = 32'h00000000;
assign filter_banks_12[116] = 32'h00000000;
assign filter_banks_12[117] = 32'h00000000;
assign filter_banks_12[118] = 32'h00000000;
assign filter_banks_12[119] = 32'h00000000;
assign filter_banks_12[120] = 32'h00000000;
assign filter_banks_12[121] = 32'h00000000;
assign filter_banks_12[122] = 32'h00000000;
assign filter_banks_12[123] = 32'h00000000;
assign filter_banks_12[124] = 32'h00000000;
assign filter_banks_12[125] = 32'h00000000;
assign filter_banks_12[126] = 32'h00000000;
assign filter_banks_12[127] = 32'h00000000;
assign filter_banks_12[128] = 32'h00000000;
assign filter_banks_12[129] = 32'h00000000;
assign filter_banks_12[130] = 32'h00000000;
assign filter_banks_12[131] = 32'h00000000;
assign filter_banks_12[132] = 32'h00000000;
assign filter_banks_12[133] = 32'h00000000;
assign filter_banks_12[134] = 32'h00000000;
assign filter_banks_12[135] = 32'h00000000;
assign filter_banks_12[136] = 32'h00000000;
assign filter_banks_12[137] = 32'h00000000;
assign filter_banks_12[138] = 32'h00000000;
assign filter_banks_12[139] = 32'h00000000;
assign filter_banks_12[140] = 32'h00000000;
assign filter_banks_12[141] = 32'h00000000;
assign filter_banks_12[142] = 32'h00000000;
assign filter_banks_12[143] = 32'h00000000;
assign filter_banks_12[144] = 32'h00000000;
assign filter_banks_12[145] = 32'h00000000;
assign filter_banks_12[146] = 32'h00000000;
assign filter_banks_12[147] = 32'h00000000;
assign filter_banks_12[148] = 32'h00000000;
assign filter_banks_12[149] = 32'h00000000;
assign filter_banks_12[150] = 32'h00000000;
assign filter_banks_12[151] = 32'h00000000;
assign filter_banks_12[152] = 32'h00000000;
assign filter_banks_12[153] = 32'h00000000;
assign filter_banks_12[154] = 32'h00000000;
assign filter_banks_12[155] = 32'h00000000;
assign filter_banks_12[156] = 32'h00000000;
assign filter_banks_12[157] = 32'h00000000;
assign filter_banks_12[158] = 32'h00000000;
assign filter_banks_12[159] = 32'h00000000;
assign filter_banks_12[160] = 32'h00000000;
assign filter_banks_12[161] = 32'h00000000;
assign filter_banks_12[162] = 32'h00000000;
assign filter_banks_12[163] = 32'h00000000;
assign filter_banks_12[164] = 32'h00000000;
assign filter_banks_12[165] = 32'h00000000;
assign filter_banks_12[166] = 32'h00000000;
assign filter_banks_12[167] = 32'h00000000;
assign filter_banks_12[168] = 32'h00000000;
assign filter_banks_12[169] = 32'h00000000;
assign filter_banks_12[170] = 32'h00000000;
assign filter_banks_12[171] = 32'h00000000;
assign filter_banks_12[172] = 32'h00000000;
assign filter_banks_12[173] = 32'h00000000;
assign filter_banks_12[174] = 32'h00000000;
assign filter_banks_12[175] = 32'h00000000;
assign filter_banks_12[176] = 32'h00000000;
assign filter_banks_12[177] = 32'h00000000;
assign filter_banks_12[178] = 32'h00000000;
assign filter_banks_12[179] = 32'h00000000;
assign filter_banks_12[180] = 32'h00000000;
assign filter_banks_12[181] = 32'h00000000;
assign filter_banks_12[182] = 32'h00000000;
assign filter_banks_12[183] = 32'h00000000;
assign filter_banks_12[184] = 32'h00000000;
assign filter_banks_12[185] = 32'h00000000;
assign filter_banks_12[186] = 32'h00000000;
assign filter_banks_12[187] = 32'h00000000;
assign filter_banks_12[188] = 32'h00000000;
assign filter_banks_12[189] = 32'h00000000;
assign filter_banks_12[190] = 32'h00000000;
assign filter_banks_12[191] = 32'h00000000;
assign filter_banks_12[192] = 32'h00000000;
assign filter_banks_12[193] = 32'h00000000;
assign filter_banks_12[194] = 32'h00000000;
assign filter_banks_12[195] = 32'h00000000;
assign filter_banks_12[196] = 32'h00000000;
assign filter_banks_12[197] = 32'h00000000;
assign filter_banks_12[198] = 32'h00000000;
assign filter_banks_12[199] = 32'h00000000;
assign filter_banks_12[200] = 32'h00000000;
assign filter_banks_12[201] = 32'h00000000;
assign filter_banks_12[202] = 32'h00000000;
assign filter_banks_12[203] = 32'h00000000;
assign filter_banks_12[204] = 32'h00000000;
assign filter_banks_12[205] = 32'h00000000;
assign filter_banks_12[206] = 32'h00000000;
assign filter_banks_12[207] = 32'h00000000;
assign filter_banks_12[208] = 32'h00000000;
assign filter_banks_12[209] = 32'h00000000;
assign filter_banks_12[210] = 32'h00000000;
assign filter_banks_12[211] = 32'h00000000;
assign filter_banks_12[212] = 32'h00000000;
assign filter_banks_12[213] = 32'h00000000;
assign filter_banks_12[214] = 32'h00000000;
assign filter_banks_12[215] = 32'h00000000;
assign filter_banks_12[216] = 32'h00000000;
assign filter_banks_12[217] = 32'h00000000;
assign filter_banks_12[218] = 32'h00000000;
assign filter_banks_12[219] = 32'h00000000;
assign filter_banks_12[220] = 32'h00000000;
assign filter_banks_12[221] = 32'h00000000;
assign filter_banks_12[222] = 32'h00000000;
assign filter_banks_12[223] = 32'h00000000;
assign filter_banks_12[224] = 32'h00000000;
assign filter_banks_12[225] = 32'h00000000;
assign filter_banks_12[226] = 32'h00000000;
assign filter_banks_12[227] = 32'h00000000;
assign filter_banks_12[228] = 32'h00000000;
assign filter_banks_12[229] = 32'h00000000;
assign filter_banks_12[230] = 32'h00000000;
assign filter_banks_12[231] = 32'h00000000;
assign filter_banks_12[232] = 32'h00000000;
assign filter_banks_12[233] = 32'h00000000;
assign filter_banks_12[234] = 32'h00000000;
assign filter_banks_12[235] = 32'h00000000;
assign filter_banks_12[236] = 32'h00000000;
assign filter_banks_12[237] = 32'h00000000;
assign filter_banks_12[238] = 32'h00000000;
assign filter_banks_12[239] = 32'h00000000;
assign filter_banks_12[240] = 32'h00000000;
assign filter_banks_12[241] = 32'h00000000;
assign filter_banks_12[242] = 32'h00000000;
assign filter_banks_12[243] = 32'h00000000;
assign filter_banks_12[244] = 32'h00000000;
assign filter_banks_12[245] = 32'h00000000;
assign filter_banks_12[246] = 32'h00000000;
assign filter_banks_12[247] = 32'h00000000;
assign filter_banks_12[248] = 32'h00000000;
assign filter_banks_12[249] = 32'h00000000;
assign filter_banks_12[250] = 32'h00000000;
assign filter_banks_12[251] = 32'h00000000;
assign filter_banks_12[252] = 32'h00000000;
assign filter_banks_12[253] = 32'h00000000;
assign filter_banks_12[254] = 32'h00000000;
assign filter_banks_12[255] = 32'h00000000;
assign filter_banks_12[256] = 32'h00000000;
assign filter_banks_13[0] = 32'h00000000;
assign filter_banks_13[1] = 32'h00000000;
assign filter_banks_13[2] = 32'h00000000;
assign filter_banks_13[3] = 32'h00000000;
assign filter_banks_13[4] = 32'h00000000;
assign filter_banks_13[5] = 32'h00000000;
assign filter_banks_13[6] = 32'h00000000;
assign filter_banks_13[7] = 32'h00000000;
assign filter_banks_13[8] = 32'h00000000;
assign filter_banks_13[9] = 32'h00000000;
assign filter_banks_13[10] = 32'h00000000;
assign filter_banks_13[11] = 32'h00000000;
assign filter_banks_13[12] = 32'h00000000;
assign filter_banks_13[13] = 32'h00000000;
assign filter_banks_13[14] = 32'h00000000;
assign filter_banks_13[15] = 32'h00000000;
assign filter_banks_13[16] = 32'h00000000;
assign filter_banks_13[17] = 32'h00000000;
assign filter_banks_13[18] = 32'h00000000;
assign filter_banks_13[19] = 32'h00000000;
assign filter_banks_13[20] = 32'h00000000;
assign filter_banks_13[21] = 32'h00000000;
assign filter_banks_13[22] = 32'h00000000;
assign filter_banks_13[23] = 32'h00000000;
assign filter_banks_13[24] = 32'h00000000;
assign filter_banks_13[25] = 32'h00000000;
assign filter_banks_13[26] = 32'h00000000;
assign filter_banks_13[27] = 32'h00000000;
assign filter_banks_13[28] = 32'h00000000;
assign filter_banks_13[29] = 32'h00000000;
assign filter_banks_13[30] = 32'h00000000;
assign filter_banks_13[31] = 32'h00000000;
assign filter_banks_13[32] = 32'h00000000;
assign filter_banks_13[33] = 32'h00000000;
assign filter_banks_13[34] = 32'h00000000;
assign filter_banks_13[35] = 32'h00000000;
assign filter_banks_13[36] = 32'h00000000;
assign filter_banks_13[37] = 32'h00000000;
assign filter_banks_13[38] = 32'h00000000;
assign filter_banks_13[39] = 32'h00000000;
assign filter_banks_13[40] = 32'h00000000;
assign filter_banks_13[41] = 32'h00000000;
assign filter_banks_13[42] = 32'h00000000;
assign filter_banks_13[43] = 32'h00000000;
assign filter_banks_13[44] = 32'h00000000;
assign filter_banks_13[45] = 32'h00000000;
assign filter_banks_13[46] = 32'h00000000;
assign filter_banks_13[47] = 32'h3e124925;
assign filter_banks_13[48] = 32'h3e924925;
assign filter_banks_13[49] = 32'h3edb6db7;
assign filter_banks_13[50] = 32'h3f124925;
assign filter_banks_13[51] = 32'h3f36db6e;
assign filter_banks_13[52] = 32'h3f5b6db7;
assign filter_banks_13[53] = 32'h3f800000;
assign filter_banks_13[54] = 32'h3f5b6db7;
assign filter_banks_13[55] = 32'h3f36db6e;
assign filter_banks_13[56] = 32'h3f124925;
assign filter_banks_13[57] = 32'h3edb6db7;
assign filter_banks_13[58] = 32'h3e924925;
assign filter_banks_13[59] = 32'h3e124925;
assign filter_banks_13[60] = 32'h00000000;
assign filter_banks_13[61] = 32'h00000000;
assign filter_banks_13[62] = 32'h00000000;
assign filter_banks_13[63] = 32'h00000000;
assign filter_banks_13[64] = 32'h00000000;
assign filter_banks_13[65] = 32'h00000000;
assign filter_banks_13[66] = 32'h00000000;
assign filter_banks_13[67] = 32'h00000000;
assign filter_banks_13[68] = 32'h00000000;
assign filter_banks_13[69] = 32'h00000000;
assign filter_banks_13[70] = 32'h00000000;
assign filter_banks_13[71] = 32'h00000000;
assign filter_banks_13[72] = 32'h00000000;
assign filter_banks_13[73] = 32'h00000000;
assign filter_banks_13[74] = 32'h00000000;
assign filter_banks_13[75] = 32'h00000000;
assign filter_banks_13[76] = 32'h00000000;
assign filter_banks_13[77] = 32'h00000000;
assign filter_banks_13[78] = 32'h00000000;
assign filter_banks_13[79] = 32'h00000000;
assign filter_banks_13[80] = 32'h00000000;
assign filter_banks_13[81] = 32'h00000000;
assign filter_banks_13[82] = 32'h00000000;
assign filter_banks_13[83] = 32'h00000000;
assign filter_banks_13[84] = 32'h00000000;
assign filter_banks_13[85] = 32'h00000000;
assign filter_banks_13[86] = 32'h00000000;
assign filter_banks_13[87] = 32'h00000000;
assign filter_banks_13[88] = 32'h00000000;
assign filter_banks_13[89] = 32'h00000000;
assign filter_banks_13[90] = 32'h00000000;
assign filter_banks_13[91] = 32'h00000000;
assign filter_banks_13[92] = 32'h00000000;
assign filter_banks_13[93] = 32'h00000000;
assign filter_banks_13[94] = 32'h00000000;
assign filter_banks_13[95] = 32'h00000000;
assign filter_banks_13[96] = 32'h00000000;
assign filter_banks_13[97] = 32'h00000000;
assign filter_banks_13[98] = 32'h00000000;
assign filter_banks_13[99] = 32'h00000000;
assign filter_banks_13[100] = 32'h00000000;
assign filter_banks_13[101] = 32'h00000000;
assign filter_banks_13[102] = 32'h00000000;
assign filter_banks_13[103] = 32'h00000000;
assign filter_banks_13[104] = 32'h00000000;
assign filter_banks_13[105] = 32'h00000000;
assign filter_banks_13[106] = 32'h00000000;
assign filter_banks_13[107] = 32'h00000000;
assign filter_banks_13[108] = 32'h00000000;
assign filter_banks_13[109] = 32'h00000000;
assign filter_banks_13[110] = 32'h00000000;
assign filter_banks_13[111] = 32'h00000000;
assign filter_banks_13[112] = 32'h00000000;
assign filter_banks_13[113] = 32'h00000000;
assign filter_banks_13[114] = 32'h00000000;
assign filter_banks_13[115] = 32'h00000000;
assign filter_banks_13[116] = 32'h00000000;
assign filter_banks_13[117] = 32'h00000000;
assign filter_banks_13[118] = 32'h00000000;
assign filter_banks_13[119] = 32'h00000000;
assign filter_banks_13[120] = 32'h00000000;
assign filter_banks_13[121] = 32'h00000000;
assign filter_banks_13[122] = 32'h00000000;
assign filter_banks_13[123] = 32'h00000000;
assign filter_banks_13[124] = 32'h00000000;
assign filter_banks_13[125] = 32'h00000000;
assign filter_banks_13[126] = 32'h00000000;
assign filter_banks_13[127] = 32'h00000000;
assign filter_banks_13[128] = 32'h00000000;
assign filter_banks_13[129] = 32'h00000000;
assign filter_banks_13[130] = 32'h00000000;
assign filter_banks_13[131] = 32'h00000000;
assign filter_banks_13[132] = 32'h00000000;
assign filter_banks_13[133] = 32'h00000000;
assign filter_banks_13[134] = 32'h00000000;
assign filter_banks_13[135] = 32'h00000000;
assign filter_banks_13[136] = 32'h00000000;
assign filter_banks_13[137] = 32'h00000000;
assign filter_banks_13[138] = 32'h00000000;
assign filter_banks_13[139] = 32'h00000000;
assign filter_banks_13[140] = 32'h00000000;
assign filter_banks_13[141] = 32'h00000000;
assign filter_banks_13[142] = 32'h00000000;
assign filter_banks_13[143] = 32'h00000000;
assign filter_banks_13[144] = 32'h00000000;
assign filter_banks_13[145] = 32'h00000000;
assign filter_banks_13[146] = 32'h00000000;
assign filter_banks_13[147] = 32'h00000000;
assign filter_banks_13[148] = 32'h00000000;
assign filter_banks_13[149] = 32'h00000000;
assign filter_banks_13[150] = 32'h00000000;
assign filter_banks_13[151] = 32'h00000000;
assign filter_banks_13[152] = 32'h00000000;
assign filter_banks_13[153] = 32'h00000000;
assign filter_banks_13[154] = 32'h00000000;
assign filter_banks_13[155] = 32'h00000000;
assign filter_banks_13[156] = 32'h00000000;
assign filter_banks_13[157] = 32'h00000000;
assign filter_banks_13[158] = 32'h00000000;
assign filter_banks_13[159] = 32'h00000000;
assign filter_banks_13[160] = 32'h00000000;
assign filter_banks_13[161] = 32'h00000000;
assign filter_banks_13[162] = 32'h00000000;
assign filter_banks_13[163] = 32'h00000000;
assign filter_banks_13[164] = 32'h00000000;
assign filter_banks_13[165] = 32'h00000000;
assign filter_banks_13[166] = 32'h00000000;
assign filter_banks_13[167] = 32'h00000000;
assign filter_banks_13[168] = 32'h00000000;
assign filter_banks_13[169] = 32'h00000000;
assign filter_banks_13[170] = 32'h00000000;
assign filter_banks_13[171] = 32'h00000000;
assign filter_banks_13[172] = 32'h00000000;
assign filter_banks_13[173] = 32'h00000000;
assign filter_banks_13[174] = 32'h00000000;
assign filter_banks_13[175] = 32'h00000000;
assign filter_banks_13[176] = 32'h00000000;
assign filter_banks_13[177] = 32'h00000000;
assign filter_banks_13[178] = 32'h00000000;
assign filter_banks_13[179] = 32'h00000000;
assign filter_banks_13[180] = 32'h00000000;
assign filter_banks_13[181] = 32'h00000000;
assign filter_banks_13[182] = 32'h00000000;
assign filter_banks_13[183] = 32'h00000000;
assign filter_banks_13[184] = 32'h00000000;
assign filter_banks_13[185] = 32'h00000000;
assign filter_banks_13[186] = 32'h00000000;
assign filter_banks_13[187] = 32'h00000000;
assign filter_banks_13[188] = 32'h00000000;
assign filter_banks_13[189] = 32'h00000000;
assign filter_banks_13[190] = 32'h00000000;
assign filter_banks_13[191] = 32'h00000000;
assign filter_banks_13[192] = 32'h00000000;
assign filter_banks_13[193] = 32'h00000000;
assign filter_banks_13[194] = 32'h00000000;
assign filter_banks_13[195] = 32'h00000000;
assign filter_banks_13[196] = 32'h00000000;
assign filter_banks_13[197] = 32'h00000000;
assign filter_banks_13[198] = 32'h00000000;
assign filter_banks_13[199] = 32'h00000000;
assign filter_banks_13[200] = 32'h00000000;
assign filter_banks_13[201] = 32'h00000000;
assign filter_banks_13[202] = 32'h00000000;
assign filter_banks_13[203] = 32'h00000000;
assign filter_banks_13[204] = 32'h00000000;
assign filter_banks_13[205] = 32'h00000000;
assign filter_banks_13[206] = 32'h00000000;
assign filter_banks_13[207] = 32'h00000000;
assign filter_banks_13[208] = 32'h00000000;
assign filter_banks_13[209] = 32'h00000000;
assign filter_banks_13[210] = 32'h00000000;
assign filter_banks_13[211] = 32'h00000000;
assign filter_banks_13[212] = 32'h00000000;
assign filter_banks_13[213] = 32'h00000000;
assign filter_banks_13[214] = 32'h00000000;
assign filter_banks_13[215] = 32'h00000000;
assign filter_banks_13[216] = 32'h00000000;
assign filter_banks_13[217] = 32'h00000000;
assign filter_banks_13[218] = 32'h00000000;
assign filter_banks_13[219] = 32'h00000000;
assign filter_banks_13[220] = 32'h00000000;
assign filter_banks_13[221] = 32'h00000000;
assign filter_banks_13[222] = 32'h00000000;
assign filter_banks_13[223] = 32'h00000000;
assign filter_banks_13[224] = 32'h00000000;
assign filter_banks_13[225] = 32'h00000000;
assign filter_banks_13[226] = 32'h00000000;
assign filter_banks_13[227] = 32'h00000000;
assign filter_banks_13[228] = 32'h00000000;
assign filter_banks_13[229] = 32'h00000000;
assign filter_banks_13[230] = 32'h00000000;
assign filter_banks_13[231] = 32'h00000000;
assign filter_banks_13[232] = 32'h00000000;
assign filter_banks_13[233] = 32'h00000000;
assign filter_banks_13[234] = 32'h00000000;
assign filter_banks_13[235] = 32'h00000000;
assign filter_banks_13[236] = 32'h00000000;
assign filter_banks_13[237] = 32'h00000000;
assign filter_banks_13[238] = 32'h00000000;
assign filter_banks_13[239] = 32'h00000000;
assign filter_banks_13[240] = 32'h00000000;
assign filter_banks_13[241] = 32'h00000000;
assign filter_banks_13[242] = 32'h00000000;
assign filter_banks_13[243] = 32'h00000000;
assign filter_banks_13[244] = 32'h00000000;
assign filter_banks_13[245] = 32'h00000000;
assign filter_banks_13[246] = 32'h00000000;
assign filter_banks_13[247] = 32'h00000000;
assign filter_banks_13[248] = 32'h00000000;
assign filter_banks_13[249] = 32'h00000000;
assign filter_banks_13[250] = 32'h00000000;
assign filter_banks_13[251] = 32'h00000000;
assign filter_banks_13[252] = 32'h00000000;
assign filter_banks_13[253] = 32'h00000000;
assign filter_banks_13[254] = 32'h00000000;
assign filter_banks_13[255] = 32'h00000000;
assign filter_banks_13[256] = 32'h00000000;
assign filter_banks_14[0] = 32'h00000000;
assign filter_banks_14[1] = 32'h00000000;
assign filter_banks_14[2] = 32'h00000000;
assign filter_banks_14[3] = 32'h00000000;
assign filter_banks_14[4] = 32'h00000000;
assign filter_banks_14[5] = 32'h00000000;
assign filter_banks_14[6] = 32'h00000000;
assign filter_banks_14[7] = 32'h00000000;
assign filter_banks_14[8] = 32'h00000000;
assign filter_banks_14[9] = 32'h00000000;
assign filter_banks_14[10] = 32'h00000000;
assign filter_banks_14[11] = 32'h00000000;
assign filter_banks_14[12] = 32'h00000000;
assign filter_banks_14[13] = 32'h00000000;
assign filter_banks_14[14] = 32'h00000000;
assign filter_banks_14[15] = 32'h00000000;
assign filter_banks_14[16] = 32'h00000000;
assign filter_banks_14[17] = 32'h00000000;
assign filter_banks_14[18] = 32'h00000000;
assign filter_banks_14[19] = 32'h00000000;
assign filter_banks_14[20] = 32'h00000000;
assign filter_banks_14[21] = 32'h00000000;
assign filter_banks_14[22] = 32'h00000000;
assign filter_banks_14[23] = 32'h00000000;
assign filter_banks_14[24] = 32'h00000000;
assign filter_banks_14[25] = 32'h00000000;
assign filter_banks_14[26] = 32'h00000000;
assign filter_banks_14[27] = 32'h00000000;
assign filter_banks_14[28] = 32'h00000000;
assign filter_banks_14[29] = 32'h00000000;
assign filter_banks_14[30] = 32'h00000000;
assign filter_banks_14[31] = 32'h00000000;
assign filter_banks_14[32] = 32'h00000000;
assign filter_banks_14[33] = 32'h00000000;
assign filter_banks_14[34] = 32'h00000000;
assign filter_banks_14[35] = 32'h00000000;
assign filter_banks_14[36] = 32'h00000000;
assign filter_banks_14[37] = 32'h00000000;
assign filter_banks_14[38] = 32'h00000000;
assign filter_banks_14[39] = 32'h00000000;
assign filter_banks_14[40] = 32'h00000000;
assign filter_banks_14[41] = 32'h00000000;
assign filter_banks_14[42] = 32'h00000000;
assign filter_banks_14[43] = 32'h00000000;
assign filter_banks_14[44] = 32'h00000000;
assign filter_banks_14[45] = 32'h00000000;
assign filter_banks_14[46] = 32'h00000000;
assign filter_banks_14[47] = 32'h00000000;
assign filter_banks_14[48] = 32'h00000000;
assign filter_banks_14[49] = 32'h00000000;
assign filter_banks_14[50] = 32'h00000000;
assign filter_banks_14[51] = 32'h00000000;
assign filter_banks_14[52] = 32'h00000000;
assign filter_banks_14[53] = 32'h00000000;
assign filter_banks_14[54] = 32'h3e124925;
assign filter_banks_14[55] = 32'h3e924925;
assign filter_banks_14[56] = 32'h3edb6db7;
assign filter_banks_14[57] = 32'h3f124925;
assign filter_banks_14[58] = 32'h3f36db6e;
assign filter_banks_14[59] = 32'h3f5b6db7;
assign filter_banks_14[60] = 32'h3f800000;
assign filter_banks_14[61] = 32'h3f600000;
assign filter_banks_14[62] = 32'h3f400000;
assign filter_banks_14[63] = 32'h3f200000;
assign filter_banks_14[64] = 32'h3f000000;
assign filter_banks_14[65] = 32'h3ec00000;
assign filter_banks_14[66] = 32'h3e800000;
assign filter_banks_14[67] = 32'h3e000000;
assign filter_banks_14[68] = 32'h00000000;
assign filter_banks_14[69] = 32'h00000000;
assign filter_banks_14[70] = 32'h00000000;
assign filter_banks_14[71] = 32'h00000000;
assign filter_banks_14[72] = 32'h00000000;
assign filter_banks_14[73] = 32'h00000000;
assign filter_banks_14[74] = 32'h00000000;
assign filter_banks_14[75] = 32'h00000000;
assign filter_banks_14[76] = 32'h00000000;
assign filter_banks_14[77] = 32'h00000000;
assign filter_banks_14[78] = 32'h00000000;
assign filter_banks_14[79] = 32'h00000000;
assign filter_banks_14[80] = 32'h00000000;
assign filter_banks_14[81] = 32'h00000000;
assign filter_banks_14[82] = 32'h00000000;
assign filter_banks_14[83] = 32'h00000000;
assign filter_banks_14[84] = 32'h00000000;
assign filter_banks_14[85] = 32'h00000000;
assign filter_banks_14[86] = 32'h00000000;
assign filter_banks_14[87] = 32'h00000000;
assign filter_banks_14[88] = 32'h00000000;
assign filter_banks_14[89] = 32'h00000000;
assign filter_banks_14[90] = 32'h00000000;
assign filter_banks_14[91] = 32'h00000000;
assign filter_banks_14[92] = 32'h00000000;
assign filter_banks_14[93] = 32'h00000000;
assign filter_banks_14[94] = 32'h00000000;
assign filter_banks_14[95] = 32'h00000000;
assign filter_banks_14[96] = 32'h00000000;
assign filter_banks_14[97] = 32'h00000000;
assign filter_banks_14[98] = 32'h00000000;
assign filter_banks_14[99] = 32'h00000000;
assign filter_banks_14[100] = 32'h00000000;
assign filter_banks_14[101] = 32'h00000000;
assign filter_banks_14[102] = 32'h00000000;
assign filter_banks_14[103] = 32'h00000000;
assign filter_banks_14[104] = 32'h00000000;
assign filter_banks_14[105] = 32'h00000000;
assign filter_banks_14[106] = 32'h00000000;
assign filter_banks_14[107] = 32'h00000000;
assign filter_banks_14[108] = 32'h00000000;
assign filter_banks_14[109] = 32'h00000000;
assign filter_banks_14[110] = 32'h00000000;
assign filter_banks_14[111] = 32'h00000000;
assign filter_banks_14[112] = 32'h00000000;
assign filter_banks_14[113] = 32'h00000000;
assign filter_banks_14[114] = 32'h00000000;
assign filter_banks_14[115] = 32'h00000000;
assign filter_banks_14[116] = 32'h00000000;
assign filter_banks_14[117] = 32'h00000000;
assign filter_banks_14[118] = 32'h00000000;
assign filter_banks_14[119] = 32'h00000000;
assign filter_banks_14[120] = 32'h00000000;
assign filter_banks_14[121] = 32'h00000000;
assign filter_banks_14[122] = 32'h00000000;
assign filter_banks_14[123] = 32'h00000000;
assign filter_banks_14[124] = 32'h00000000;
assign filter_banks_14[125] = 32'h00000000;
assign filter_banks_14[126] = 32'h00000000;
assign filter_banks_14[127] = 32'h00000000;
assign filter_banks_14[128] = 32'h00000000;
assign filter_banks_14[129] = 32'h00000000;
assign filter_banks_14[130] = 32'h00000000;
assign filter_banks_14[131] = 32'h00000000;
assign filter_banks_14[132] = 32'h00000000;
assign filter_banks_14[133] = 32'h00000000;
assign filter_banks_14[134] = 32'h00000000;
assign filter_banks_14[135] = 32'h00000000;
assign filter_banks_14[136] = 32'h00000000;
assign filter_banks_14[137] = 32'h00000000;
assign filter_banks_14[138] = 32'h00000000;
assign filter_banks_14[139] = 32'h00000000;
assign filter_banks_14[140] = 32'h00000000;
assign filter_banks_14[141] = 32'h00000000;
assign filter_banks_14[142] = 32'h00000000;
assign filter_banks_14[143] = 32'h00000000;
assign filter_banks_14[144] = 32'h00000000;
assign filter_banks_14[145] = 32'h00000000;
assign filter_banks_14[146] = 32'h00000000;
assign filter_banks_14[147] = 32'h00000000;
assign filter_banks_14[148] = 32'h00000000;
assign filter_banks_14[149] = 32'h00000000;
assign filter_banks_14[150] = 32'h00000000;
assign filter_banks_14[151] = 32'h00000000;
assign filter_banks_14[152] = 32'h00000000;
assign filter_banks_14[153] = 32'h00000000;
assign filter_banks_14[154] = 32'h00000000;
assign filter_banks_14[155] = 32'h00000000;
assign filter_banks_14[156] = 32'h00000000;
assign filter_banks_14[157] = 32'h00000000;
assign filter_banks_14[158] = 32'h00000000;
assign filter_banks_14[159] = 32'h00000000;
assign filter_banks_14[160] = 32'h00000000;
assign filter_banks_14[161] = 32'h00000000;
assign filter_banks_14[162] = 32'h00000000;
assign filter_banks_14[163] = 32'h00000000;
assign filter_banks_14[164] = 32'h00000000;
assign filter_banks_14[165] = 32'h00000000;
assign filter_banks_14[166] = 32'h00000000;
assign filter_banks_14[167] = 32'h00000000;
assign filter_banks_14[168] = 32'h00000000;
assign filter_banks_14[169] = 32'h00000000;
assign filter_banks_14[170] = 32'h00000000;
assign filter_banks_14[171] = 32'h00000000;
assign filter_banks_14[172] = 32'h00000000;
assign filter_banks_14[173] = 32'h00000000;
assign filter_banks_14[174] = 32'h00000000;
assign filter_banks_14[175] = 32'h00000000;
assign filter_banks_14[176] = 32'h00000000;
assign filter_banks_14[177] = 32'h00000000;
assign filter_banks_14[178] = 32'h00000000;
assign filter_banks_14[179] = 32'h00000000;
assign filter_banks_14[180] = 32'h00000000;
assign filter_banks_14[181] = 32'h00000000;
assign filter_banks_14[182] = 32'h00000000;
assign filter_banks_14[183] = 32'h00000000;
assign filter_banks_14[184] = 32'h00000000;
assign filter_banks_14[185] = 32'h00000000;
assign filter_banks_14[186] = 32'h00000000;
assign filter_banks_14[187] = 32'h00000000;
assign filter_banks_14[188] = 32'h00000000;
assign filter_banks_14[189] = 32'h00000000;
assign filter_banks_14[190] = 32'h00000000;
assign filter_banks_14[191] = 32'h00000000;
assign filter_banks_14[192] = 32'h00000000;
assign filter_banks_14[193] = 32'h00000000;
assign filter_banks_14[194] = 32'h00000000;
assign filter_banks_14[195] = 32'h00000000;
assign filter_banks_14[196] = 32'h00000000;
assign filter_banks_14[197] = 32'h00000000;
assign filter_banks_14[198] = 32'h00000000;
assign filter_banks_14[199] = 32'h00000000;
assign filter_banks_14[200] = 32'h00000000;
assign filter_banks_14[201] = 32'h00000000;
assign filter_banks_14[202] = 32'h00000000;
assign filter_banks_14[203] = 32'h00000000;
assign filter_banks_14[204] = 32'h00000000;
assign filter_banks_14[205] = 32'h00000000;
assign filter_banks_14[206] = 32'h00000000;
assign filter_banks_14[207] = 32'h00000000;
assign filter_banks_14[208] = 32'h00000000;
assign filter_banks_14[209] = 32'h00000000;
assign filter_banks_14[210] = 32'h00000000;
assign filter_banks_14[211] = 32'h00000000;
assign filter_banks_14[212] = 32'h00000000;
assign filter_banks_14[213] = 32'h00000000;
assign filter_banks_14[214] = 32'h00000000;
assign filter_banks_14[215] = 32'h00000000;
assign filter_banks_14[216] = 32'h00000000;
assign filter_banks_14[217] = 32'h00000000;
assign filter_banks_14[218] = 32'h00000000;
assign filter_banks_14[219] = 32'h00000000;
assign filter_banks_14[220] = 32'h00000000;
assign filter_banks_14[221] = 32'h00000000;
assign filter_banks_14[222] = 32'h00000000;
assign filter_banks_14[223] = 32'h00000000;
assign filter_banks_14[224] = 32'h00000000;
assign filter_banks_14[225] = 32'h00000000;
assign filter_banks_14[226] = 32'h00000000;
assign filter_banks_14[227] = 32'h00000000;
assign filter_banks_14[228] = 32'h00000000;
assign filter_banks_14[229] = 32'h00000000;
assign filter_banks_14[230] = 32'h00000000;
assign filter_banks_14[231] = 32'h00000000;
assign filter_banks_14[232] = 32'h00000000;
assign filter_banks_14[233] = 32'h00000000;
assign filter_banks_14[234] = 32'h00000000;
assign filter_banks_14[235] = 32'h00000000;
assign filter_banks_14[236] = 32'h00000000;
assign filter_banks_14[237] = 32'h00000000;
assign filter_banks_14[238] = 32'h00000000;
assign filter_banks_14[239] = 32'h00000000;
assign filter_banks_14[240] = 32'h00000000;
assign filter_banks_14[241] = 32'h00000000;
assign filter_banks_14[242] = 32'h00000000;
assign filter_banks_14[243] = 32'h00000000;
assign filter_banks_14[244] = 32'h00000000;
assign filter_banks_14[245] = 32'h00000000;
assign filter_banks_14[246] = 32'h00000000;
assign filter_banks_14[247] = 32'h00000000;
assign filter_banks_14[248] = 32'h00000000;
assign filter_banks_14[249] = 32'h00000000;
assign filter_banks_14[250] = 32'h00000000;
assign filter_banks_14[251] = 32'h00000000;
assign filter_banks_14[252] = 32'h00000000;
assign filter_banks_14[253] = 32'h00000000;
assign filter_banks_14[254] = 32'h00000000;
assign filter_banks_14[255] = 32'h00000000;
assign filter_banks_14[256] = 32'h00000000;
assign filter_banks_15[0] = 32'h00000000;
assign filter_banks_15[1] = 32'h00000000;
assign filter_banks_15[2] = 32'h00000000;
assign filter_banks_15[3] = 32'h00000000;
assign filter_banks_15[4] = 32'h00000000;
assign filter_banks_15[5] = 32'h00000000;
assign filter_banks_15[6] = 32'h00000000;
assign filter_banks_15[7] = 32'h00000000;
assign filter_banks_15[8] = 32'h00000000;
assign filter_banks_15[9] = 32'h00000000;
assign filter_banks_15[10] = 32'h00000000;
assign filter_banks_15[11] = 32'h00000000;
assign filter_banks_15[12] = 32'h00000000;
assign filter_banks_15[13] = 32'h00000000;
assign filter_banks_15[14] = 32'h00000000;
assign filter_banks_15[15] = 32'h00000000;
assign filter_banks_15[16] = 32'h00000000;
assign filter_banks_15[17] = 32'h00000000;
assign filter_banks_15[18] = 32'h00000000;
assign filter_banks_15[19] = 32'h00000000;
assign filter_banks_15[20] = 32'h00000000;
assign filter_banks_15[21] = 32'h00000000;
assign filter_banks_15[22] = 32'h00000000;
assign filter_banks_15[23] = 32'h00000000;
assign filter_banks_15[24] = 32'h00000000;
assign filter_banks_15[25] = 32'h00000000;
assign filter_banks_15[26] = 32'h00000000;
assign filter_banks_15[27] = 32'h00000000;
assign filter_banks_15[28] = 32'h00000000;
assign filter_banks_15[29] = 32'h00000000;
assign filter_banks_15[30] = 32'h00000000;
assign filter_banks_15[31] = 32'h00000000;
assign filter_banks_15[32] = 32'h00000000;
assign filter_banks_15[33] = 32'h00000000;
assign filter_banks_15[34] = 32'h00000000;
assign filter_banks_15[35] = 32'h00000000;
assign filter_banks_15[36] = 32'h00000000;
assign filter_banks_15[37] = 32'h00000000;
assign filter_banks_15[38] = 32'h00000000;
assign filter_banks_15[39] = 32'h00000000;
assign filter_banks_15[40] = 32'h00000000;
assign filter_banks_15[41] = 32'h00000000;
assign filter_banks_15[42] = 32'h00000000;
assign filter_banks_15[43] = 32'h00000000;
assign filter_banks_15[44] = 32'h00000000;
assign filter_banks_15[45] = 32'h00000000;
assign filter_banks_15[46] = 32'h00000000;
assign filter_banks_15[47] = 32'h00000000;
assign filter_banks_15[48] = 32'h00000000;
assign filter_banks_15[49] = 32'h00000000;
assign filter_banks_15[50] = 32'h00000000;
assign filter_banks_15[51] = 32'h00000000;
assign filter_banks_15[52] = 32'h00000000;
assign filter_banks_15[53] = 32'h00000000;
assign filter_banks_15[54] = 32'h00000000;
assign filter_banks_15[55] = 32'h00000000;
assign filter_banks_15[56] = 32'h00000000;
assign filter_banks_15[57] = 32'h00000000;
assign filter_banks_15[58] = 32'h00000000;
assign filter_banks_15[59] = 32'h00000000;
assign filter_banks_15[60] = 32'h00000000;
assign filter_banks_15[61] = 32'h3e000000;
assign filter_banks_15[62] = 32'h3e800000;
assign filter_banks_15[63] = 32'h3ec00000;
assign filter_banks_15[64] = 32'h3f000000;
assign filter_banks_15[65] = 32'h3f200000;
assign filter_banks_15[66] = 32'h3f400000;
assign filter_banks_15[67] = 32'h3f600000;
assign filter_banks_15[68] = 32'h3f800000;
assign filter_banks_15[69] = 32'h3f638e39;
assign filter_banks_15[70] = 32'h3f471c72;
assign filter_banks_15[71] = 32'h3f2aaaab;
assign filter_banks_15[72] = 32'h3f0e38e4;
assign filter_banks_15[73] = 32'h3ee38e39;
assign filter_banks_15[74] = 32'h3eaaaaab;
assign filter_banks_15[75] = 32'h3e638e39;
assign filter_banks_15[76] = 32'h3de38e39;
assign filter_banks_15[77] = 32'h00000000;
assign filter_banks_15[78] = 32'h00000000;
assign filter_banks_15[79] = 32'h00000000;
assign filter_banks_15[80] = 32'h00000000;
assign filter_banks_15[81] = 32'h00000000;
assign filter_banks_15[82] = 32'h00000000;
assign filter_banks_15[83] = 32'h00000000;
assign filter_banks_15[84] = 32'h00000000;
assign filter_banks_15[85] = 32'h00000000;
assign filter_banks_15[86] = 32'h00000000;
assign filter_banks_15[87] = 32'h00000000;
assign filter_banks_15[88] = 32'h00000000;
assign filter_banks_15[89] = 32'h00000000;
assign filter_banks_15[90] = 32'h00000000;
assign filter_banks_15[91] = 32'h00000000;
assign filter_banks_15[92] = 32'h00000000;
assign filter_banks_15[93] = 32'h00000000;
assign filter_banks_15[94] = 32'h00000000;
assign filter_banks_15[95] = 32'h00000000;
assign filter_banks_15[96] = 32'h00000000;
assign filter_banks_15[97] = 32'h00000000;
assign filter_banks_15[98] = 32'h00000000;
assign filter_banks_15[99] = 32'h00000000;
assign filter_banks_15[100] = 32'h00000000;
assign filter_banks_15[101] = 32'h00000000;
assign filter_banks_15[102] = 32'h00000000;
assign filter_banks_15[103] = 32'h00000000;
assign filter_banks_15[104] = 32'h00000000;
assign filter_banks_15[105] = 32'h00000000;
assign filter_banks_15[106] = 32'h00000000;
assign filter_banks_15[107] = 32'h00000000;
assign filter_banks_15[108] = 32'h00000000;
assign filter_banks_15[109] = 32'h00000000;
assign filter_banks_15[110] = 32'h00000000;
assign filter_banks_15[111] = 32'h00000000;
assign filter_banks_15[112] = 32'h00000000;
assign filter_banks_15[113] = 32'h00000000;
assign filter_banks_15[114] = 32'h00000000;
assign filter_banks_15[115] = 32'h00000000;
assign filter_banks_15[116] = 32'h00000000;
assign filter_banks_15[117] = 32'h00000000;
assign filter_banks_15[118] = 32'h00000000;
assign filter_banks_15[119] = 32'h00000000;
assign filter_banks_15[120] = 32'h00000000;
assign filter_banks_15[121] = 32'h00000000;
assign filter_banks_15[122] = 32'h00000000;
assign filter_banks_15[123] = 32'h00000000;
assign filter_banks_15[124] = 32'h00000000;
assign filter_banks_15[125] = 32'h00000000;
assign filter_banks_15[126] = 32'h00000000;
assign filter_banks_15[127] = 32'h00000000;
assign filter_banks_15[128] = 32'h00000000;
assign filter_banks_15[129] = 32'h00000000;
assign filter_banks_15[130] = 32'h00000000;
assign filter_banks_15[131] = 32'h00000000;
assign filter_banks_15[132] = 32'h00000000;
assign filter_banks_15[133] = 32'h00000000;
assign filter_banks_15[134] = 32'h00000000;
assign filter_banks_15[135] = 32'h00000000;
assign filter_banks_15[136] = 32'h00000000;
assign filter_banks_15[137] = 32'h00000000;
assign filter_banks_15[138] = 32'h00000000;
assign filter_banks_15[139] = 32'h00000000;
assign filter_banks_15[140] = 32'h00000000;
assign filter_banks_15[141] = 32'h00000000;
assign filter_banks_15[142] = 32'h00000000;
assign filter_banks_15[143] = 32'h00000000;
assign filter_banks_15[144] = 32'h00000000;
assign filter_banks_15[145] = 32'h00000000;
assign filter_banks_15[146] = 32'h00000000;
assign filter_banks_15[147] = 32'h00000000;
assign filter_banks_15[148] = 32'h00000000;
assign filter_banks_15[149] = 32'h00000000;
assign filter_banks_15[150] = 32'h00000000;
assign filter_banks_15[151] = 32'h00000000;
assign filter_banks_15[152] = 32'h00000000;
assign filter_banks_15[153] = 32'h00000000;
assign filter_banks_15[154] = 32'h00000000;
assign filter_banks_15[155] = 32'h00000000;
assign filter_banks_15[156] = 32'h00000000;
assign filter_banks_15[157] = 32'h00000000;
assign filter_banks_15[158] = 32'h00000000;
assign filter_banks_15[159] = 32'h00000000;
assign filter_banks_15[160] = 32'h00000000;
assign filter_banks_15[161] = 32'h00000000;
assign filter_banks_15[162] = 32'h00000000;
assign filter_banks_15[163] = 32'h00000000;
assign filter_banks_15[164] = 32'h00000000;
assign filter_banks_15[165] = 32'h00000000;
assign filter_banks_15[166] = 32'h00000000;
assign filter_banks_15[167] = 32'h00000000;
assign filter_banks_15[168] = 32'h00000000;
assign filter_banks_15[169] = 32'h00000000;
assign filter_banks_15[170] = 32'h00000000;
assign filter_banks_15[171] = 32'h00000000;
assign filter_banks_15[172] = 32'h00000000;
assign filter_banks_15[173] = 32'h00000000;
assign filter_banks_15[174] = 32'h00000000;
assign filter_banks_15[175] = 32'h00000000;
assign filter_banks_15[176] = 32'h00000000;
assign filter_banks_15[177] = 32'h00000000;
assign filter_banks_15[178] = 32'h00000000;
assign filter_banks_15[179] = 32'h00000000;
assign filter_banks_15[180] = 32'h00000000;
assign filter_banks_15[181] = 32'h00000000;
assign filter_banks_15[182] = 32'h00000000;
assign filter_banks_15[183] = 32'h00000000;
assign filter_banks_15[184] = 32'h00000000;
assign filter_banks_15[185] = 32'h00000000;
assign filter_banks_15[186] = 32'h00000000;
assign filter_banks_15[187] = 32'h00000000;
assign filter_banks_15[188] = 32'h00000000;
assign filter_banks_15[189] = 32'h00000000;
assign filter_banks_15[190] = 32'h00000000;
assign filter_banks_15[191] = 32'h00000000;
assign filter_banks_15[192] = 32'h00000000;
assign filter_banks_15[193] = 32'h00000000;
assign filter_banks_15[194] = 32'h00000000;
assign filter_banks_15[195] = 32'h00000000;
assign filter_banks_15[196] = 32'h00000000;
assign filter_banks_15[197] = 32'h00000000;
assign filter_banks_15[198] = 32'h00000000;
assign filter_banks_15[199] = 32'h00000000;
assign filter_banks_15[200] = 32'h00000000;
assign filter_banks_15[201] = 32'h00000000;
assign filter_banks_15[202] = 32'h00000000;
assign filter_banks_15[203] = 32'h00000000;
assign filter_banks_15[204] = 32'h00000000;
assign filter_banks_15[205] = 32'h00000000;
assign filter_banks_15[206] = 32'h00000000;
assign filter_banks_15[207] = 32'h00000000;
assign filter_banks_15[208] = 32'h00000000;
assign filter_banks_15[209] = 32'h00000000;
assign filter_banks_15[210] = 32'h00000000;
assign filter_banks_15[211] = 32'h00000000;
assign filter_banks_15[212] = 32'h00000000;
assign filter_banks_15[213] = 32'h00000000;
assign filter_banks_15[214] = 32'h00000000;
assign filter_banks_15[215] = 32'h00000000;
assign filter_banks_15[216] = 32'h00000000;
assign filter_banks_15[217] = 32'h00000000;
assign filter_banks_15[218] = 32'h00000000;
assign filter_banks_15[219] = 32'h00000000;
assign filter_banks_15[220] = 32'h00000000;
assign filter_banks_15[221] = 32'h00000000;
assign filter_banks_15[222] = 32'h00000000;
assign filter_banks_15[223] = 32'h00000000;
assign filter_banks_15[224] = 32'h00000000;
assign filter_banks_15[225] = 32'h00000000;
assign filter_banks_15[226] = 32'h00000000;
assign filter_banks_15[227] = 32'h00000000;
assign filter_banks_15[228] = 32'h00000000;
assign filter_banks_15[229] = 32'h00000000;
assign filter_banks_15[230] = 32'h00000000;
assign filter_banks_15[231] = 32'h00000000;
assign filter_banks_15[232] = 32'h00000000;
assign filter_banks_15[233] = 32'h00000000;
assign filter_banks_15[234] = 32'h00000000;
assign filter_banks_15[235] = 32'h00000000;
assign filter_banks_15[236] = 32'h00000000;
assign filter_banks_15[237] = 32'h00000000;
assign filter_banks_15[238] = 32'h00000000;
assign filter_banks_15[239] = 32'h00000000;
assign filter_banks_15[240] = 32'h00000000;
assign filter_banks_15[241] = 32'h00000000;
assign filter_banks_15[242] = 32'h00000000;
assign filter_banks_15[243] = 32'h00000000;
assign filter_banks_15[244] = 32'h00000000;
assign filter_banks_15[245] = 32'h00000000;
assign filter_banks_15[246] = 32'h00000000;
assign filter_banks_15[247] = 32'h00000000;
assign filter_banks_15[248] = 32'h00000000;
assign filter_banks_15[249] = 32'h00000000;
assign filter_banks_15[250] = 32'h00000000;
assign filter_banks_15[251] = 32'h00000000;
assign filter_banks_15[252] = 32'h00000000;
assign filter_banks_15[253] = 32'h00000000;
assign filter_banks_15[254] = 32'h00000000;
assign filter_banks_15[255] = 32'h00000000;
assign filter_banks_15[256] = 32'h00000000;
assign filter_banks_16[0] = 32'h00000000;
assign filter_banks_16[1] = 32'h00000000;
assign filter_banks_16[2] = 32'h00000000;
assign filter_banks_16[3] = 32'h00000000;
assign filter_banks_16[4] = 32'h00000000;
assign filter_banks_16[5] = 32'h00000000;
assign filter_banks_16[6] = 32'h00000000;
assign filter_banks_16[7] = 32'h00000000;
assign filter_banks_16[8] = 32'h00000000;
assign filter_banks_16[9] = 32'h00000000;
assign filter_banks_16[10] = 32'h00000000;
assign filter_banks_16[11] = 32'h00000000;
assign filter_banks_16[12] = 32'h00000000;
assign filter_banks_16[13] = 32'h00000000;
assign filter_banks_16[14] = 32'h00000000;
assign filter_banks_16[15] = 32'h00000000;
assign filter_banks_16[16] = 32'h00000000;
assign filter_banks_16[17] = 32'h00000000;
assign filter_banks_16[18] = 32'h00000000;
assign filter_banks_16[19] = 32'h00000000;
assign filter_banks_16[20] = 32'h00000000;
assign filter_banks_16[21] = 32'h00000000;
assign filter_banks_16[22] = 32'h00000000;
assign filter_banks_16[23] = 32'h00000000;
assign filter_banks_16[24] = 32'h00000000;
assign filter_banks_16[25] = 32'h00000000;
assign filter_banks_16[26] = 32'h00000000;
assign filter_banks_16[27] = 32'h00000000;
assign filter_banks_16[28] = 32'h00000000;
assign filter_banks_16[29] = 32'h00000000;
assign filter_banks_16[30] = 32'h00000000;
assign filter_banks_16[31] = 32'h00000000;
assign filter_banks_16[32] = 32'h00000000;
assign filter_banks_16[33] = 32'h00000000;
assign filter_banks_16[34] = 32'h00000000;
assign filter_banks_16[35] = 32'h00000000;
assign filter_banks_16[36] = 32'h00000000;
assign filter_banks_16[37] = 32'h00000000;
assign filter_banks_16[38] = 32'h00000000;
assign filter_banks_16[39] = 32'h00000000;
assign filter_banks_16[40] = 32'h00000000;
assign filter_banks_16[41] = 32'h00000000;
assign filter_banks_16[42] = 32'h00000000;
assign filter_banks_16[43] = 32'h00000000;
assign filter_banks_16[44] = 32'h00000000;
assign filter_banks_16[45] = 32'h00000000;
assign filter_banks_16[46] = 32'h00000000;
assign filter_banks_16[47] = 32'h00000000;
assign filter_banks_16[48] = 32'h00000000;
assign filter_banks_16[49] = 32'h00000000;
assign filter_banks_16[50] = 32'h00000000;
assign filter_banks_16[51] = 32'h00000000;
assign filter_banks_16[52] = 32'h00000000;
assign filter_banks_16[53] = 32'h00000000;
assign filter_banks_16[54] = 32'h00000000;
assign filter_banks_16[55] = 32'h00000000;
assign filter_banks_16[56] = 32'h00000000;
assign filter_banks_16[57] = 32'h00000000;
assign filter_banks_16[58] = 32'h00000000;
assign filter_banks_16[59] = 32'h00000000;
assign filter_banks_16[60] = 32'h00000000;
assign filter_banks_16[61] = 32'h00000000;
assign filter_banks_16[62] = 32'h00000000;
assign filter_banks_16[63] = 32'h00000000;
assign filter_banks_16[64] = 32'h00000000;
assign filter_banks_16[65] = 32'h00000000;
assign filter_banks_16[66] = 32'h00000000;
assign filter_banks_16[67] = 32'h00000000;
assign filter_banks_16[68] = 32'h00000000;
assign filter_banks_16[69] = 32'h3de38e39;
assign filter_banks_16[70] = 32'h3e638e39;
assign filter_banks_16[71] = 32'h3eaaaaab;
assign filter_banks_16[72] = 32'h3ee38e39;
assign filter_banks_16[73] = 32'h3f0e38e4;
assign filter_banks_16[74] = 32'h3f2aaaab;
assign filter_banks_16[75] = 32'h3f471c72;
assign filter_banks_16[76] = 32'h3f638e39;
assign filter_banks_16[77] = 32'h3f800000;
assign filter_banks_16[78] = 32'h3f666666;
assign filter_banks_16[79] = 32'h3f4ccccd;
assign filter_banks_16[80] = 32'h3f333333;
assign filter_banks_16[81] = 32'h3f19999a;
assign filter_banks_16[82] = 32'h3f000000;
assign filter_banks_16[83] = 32'h3ecccccd;
assign filter_banks_16[84] = 32'h3e99999a;
assign filter_banks_16[85] = 32'h3e4ccccd;
assign filter_banks_16[86] = 32'h3dcccccd;
assign filter_banks_16[87] = 32'h00000000;
assign filter_banks_16[88] = 32'h00000000;
assign filter_banks_16[89] = 32'h00000000;
assign filter_banks_16[90] = 32'h00000000;
assign filter_banks_16[91] = 32'h00000000;
assign filter_banks_16[92] = 32'h00000000;
assign filter_banks_16[93] = 32'h00000000;
assign filter_banks_16[94] = 32'h00000000;
assign filter_banks_16[95] = 32'h00000000;
assign filter_banks_16[96] = 32'h00000000;
assign filter_banks_16[97] = 32'h00000000;
assign filter_banks_16[98] = 32'h00000000;
assign filter_banks_16[99] = 32'h00000000;
assign filter_banks_16[100] = 32'h00000000;
assign filter_banks_16[101] = 32'h00000000;
assign filter_banks_16[102] = 32'h00000000;
assign filter_banks_16[103] = 32'h00000000;
assign filter_banks_16[104] = 32'h00000000;
assign filter_banks_16[105] = 32'h00000000;
assign filter_banks_16[106] = 32'h00000000;
assign filter_banks_16[107] = 32'h00000000;
assign filter_banks_16[108] = 32'h00000000;
assign filter_banks_16[109] = 32'h00000000;
assign filter_banks_16[110] = 32'h00000000;
assign filter_banks_16[111] = 32'h00000000;
assign filter_banks_16[112] = 32'h00000000;
assign filter_banks_16[113] = 32'h00000000;
assign filter_banks_16[114] = 32'h00000000;
assign filter_banks_16[115] = 32'h00000000;
assign filter_banks_16[116] = 32'h00000000;
assign filter_banks_16[117] = 32'h00000000;
assign filter_banks_16[118] = 32'h00000000;
assign filter_banks_16[119] = 32'h00000000;
assign filter_banks_16[120] = 32'h00000000;
assign filter_banks_16[121] = 32'h00000000;
assign filter_banks_16[122] = 32'h00000000;
assign filter_banks_16[123] = 32'h00000000;
assign filter_banks_16[124] = 32'h00000000;
assign filter_banks_16[125] = 32'h00000000;
assign filter_banks_16[126] = 32'h00000000;
assign filter_banks_16[127] = 32'h00000000;
assign filter_banks_16[128] = 32'h00000000;
assign filter_banks_16[129] = 32'h00000000;
assign filter_banks_16[130] = 32'h00000000;
assign filter_banks_16[131] = 32'h00000000;
assign filter_banks_16[132] = 32'h00000000;
assign filter_banks_16[133] = 32'h00000000;
assign filter_banks_16[134] = 32'h00000000;
assign filter_banks_16[135] = 32'h00000000;
assign filter_banks_16[136] = 32'h00000000;
assign filter_banks_16[137] = 32'h00000000;
assign filter_banks_16[138] = 32'h00000000;
assign filter_banks_16[139] = 32'h00000000;
assign filter_banks_16[140] = 32'h00000000;
assign filter_banks_16[141] = 32'h00000000;
assign filter_banks_16[142] = 32'h00000000;
assign filter_banks_16[143] = 32'h00000000;
assign filter_banks_16[144] = 32'h00000000;
assign filter_banks_16[145] = 32'h00000000;
assign filter_banks_16[146] = 32'h00000000;
assign filter_banks_16[147] = 32'h00000000;
assign filter_banks_16[148] = 32'h00000000;
assign filter_banks_16[149] = 32'h00000000;
assign filter_banks_16[150] = 32'h00000000;
assign filter_banks_16[151] = 32'h00000000;
assign filter_banks_16[152] = 32'h00000000;
assign filter_banks_16[153] = 32'h00000000;
assign filter_banks_16[154] = 32'h00000000;
assign filter_banks_16[155] = 32'h00000000;
assign filter_banks_16[156] = 32'h00000000;
assign filter_banks_16[157] = 32'h00000000;
assign filter_banks_16[158] = 32'h00000000;
assign filter_banks_16[159] = 32'h00000000;
assign filter_banks_16[160] = 32'h00000000;
assign filter_banks_16[161] = 32'h00000000;
assign filter_banks_16[162] = 32'h00000000;
assign filter_banks_16[163] = 32'h00000000;
assign filter_banks_16[164] = 32'h00000000;
assign filter_banks_16[165] = 32'h00000000;
assign filter_banks_16[166] = 32'h00000000;
assign filter_banks_16[167] = 32'h00000000;
assign filter_banks_16[168] = 32'h00000000;
assign filter_banks_16[169] = 32'h00000000;
assign filter_banks_16[170] = 32'h00000000;
assign filter_banks_16[171] = 32'h00000000;
assign filter_banks_16[172] = 32'h00000000;
assign filter_banks_16[173] = 32'h00000000;
assign filter_banks_16[174] = 32'h00000000;
assign filter_banks_16[175] = 32'h00000000;
assign filter_banks_16[176] = 32'h00000000;
assign filter_banks_16[177] = 32'h00000000;
assign filter_banks_16[178] = 32'h00000000;
assign filter_banks_16[179] = 32'h00000000;
assign filter_banks_16[180] = 32'h00000000;
assign filter_banks_16[181] = 32'h00000000;
assign filter_banks_16[182] = 32'h00000000;
assign filter_banks_16[183] = 32'h00000000;
assign filter_banks_16[184] = 32'h00000000;
assign filter_banks_16[185] = 32'h00000000;
assign filter_banks_16[186] = 32'h00000000;
assign filter_banks_16[187] = 32'h00000000;
assign filter_banks_16[188] = 32'h00000000;
assign filter_banks_16[189] = 32'h00000000;
assign filter_banks_16[190] = 32'h00000000;
assign filter_banks_16[191] = 32'h00000000;
assign filter_banks_16[192] = 32'h00000000;
assign filter_banks_16[193] = 32'h00000000;
assign filter_banks_16[194] = 32'h00000000;
assign filter_banks_16[195] = 32'h00000000;
assign filter_banks_16[196] = 32'h00000000;
assign filter_banks_16[197] = 32'h00000000;
assign filter_banks_16[198] = 32'h00000000;
assign filter_banks_16[199] = 32'h00000000;
assign filter_banks_16[200] = 32'h00000000;
assign filter_banks_16[201] = 32'h00000000;
assign filter_banks_16[202] = 32'h00000000;
assign filter_banks_16[203] = 32'h00000000;
assign filter_banks_16[204] = 32'h00000000;
assign filter_banks_16[205] = 32'h00000000;
assign filter_banks_16[206] = 32'h00000000;
assign filter_banks_16[207] = 32'h00000000;
assign filter_banks_16[208] = 32'h00000000;
assign filter_banks_16[209] = 32'h00000000;
assign filter_banks_16[210] = 32'h00000000;
assign filter_banks_16[211] = 32'h00000000;
assign filter_banks_16[212] = 32'h00000000;
assign filter_banks_16[213] = 32'h00000000;
assign filter_banks_16[214] = 32'h00000000;
assign filter_banks_16[215] = 32'h00000000;
assign filter_banks_16[216] = 32'h00000000;
assign filter_banks_16[217] = 32'h00000000;
assign filter_banks_16[218] = 32'h00000000;
assign filter_banks_16[219] = 32'h00000000;
assign filter_banks_16[220] = 32'h00000000;
assign filter_banks_16[221] = 32'h00000000;
assign filter_banks_16[222] = 32'h00000000;
assign filter_banks_16[223] = 32'h00000000;
assign filter_banks_16[224] = 32'h00000000;
assign filter_banks_16[225] = 32'h00000000;
assign filter_banks_16[226] = 32'h00000000;
assign filter_banks_16[227] = 32'h00000000;
assign filter_banks_16[228] = 32'h00000000;
assign filter_banks_16[229] = 32'h00000000;
assign filter_banks_16[230] = 32'h00000000;
assign filter_banks_16[231] = 32'h00000000;
assign filter_banks_16[232] = 32'h00000000;
assign filter_banks_16[233] = 32'h00000000;
assign filter_banks_16[234] = 32'h00000000;
assign filter_banks_16[235] = 32'h00000000;
assign filter_banks_16[236] = 32'h00000000;
assign filter_banks_16[237] = 32'h00000000;
assign filter_banks_16[238] = 32'h00000000;
assign filter_banks_16[239] = 32'h00000000;
assign filter_banks_16[240] = 32'h00000000;
assign filter_banks_16[241] = 32'h00000000;
assign filter_banks_16[242] = 32'h00000000;
assign filter_banks_16[243] = 32'h00000000;
assign filter_banks_16[244] = 32'h00000000;
assign filter_banks_16[245] = 32'h00000000;
assign filter_banks_16[246] = 32'h00000000;
assign filter_banks_16[247] = 32'h00000000;
assign filter_banks_16[248] = 32'h00000000;
assign filter_banks_16[249] = 32'h00000000;
assign filter_banks_16[250] = 32'h00000000;
assign filter_banks_16[251] = 32'h00000000;
assign filter_banks_16[252] = 32'h00000000;
assign filter_banks_16[253] = 32'h00000000;
assign filter_banks_16[254] = 32'h00000000;
assign filter_banks_16[255] = 32'h00000000;
assign filter_banks_16[256] = 32'h00000000;
assign filter_banks_17[0] = 32'h00000000;
assign filter_banks_17[1] = 32'h00000000;
assign filter_banks_17[2] = 32'h00000000;
assign filter_banks_17[3] = 32'h00000000;
assign filter_banks_17[4] = 32'h00000000;
assign filter_banks_17[5] = 32'h00000000;
assign filter_banks_17[6] = 32'h00000000;
assign filter_banks_17[7] = 32'h00000000;
assign filter_banks_17[8] = 32'h00000000;
assign filter_banks_17[9] = 32'h00000000;
assign filter_banks_17[10] = 32'h00000000;
assign filter_banks_17[11] = 32'h00000000;
assign filter_banks_17[12] = 32'h00000000;
assign filter_banks_17[13] = 32'h00000000;
assign filter_banks_17[14] = 32'h00000000;
assign filter_banks_17[15] = 32'h00000000;
assign filter_banks_17[16] = 32'h00000000;
assign filter_banks_17[17] = 32'h00000000;
assign filter_banks_17[18] = 32'h00000000;
assign filter_banks_17[19] = 32'h00000000;
assign filter_banks_17[20] = 32'h00000000;
assign filter_banks_17[21] = 32'h00000000;
assign filter_banks_17[22] = 32'h00000000;
assign filter_banks_17[23] = 32'h00000000;
assign filter_banks_17[24] = 32'h00000000;
assign filter_banks_17[25] = 32'h00000000;
assign filter_banks_17[26] = 32'h00000000;
assign filter_banks_17[27] = 32'h00000000;
assign filter_banks_17[28] = 32'h00000000;
assign filter_banks_17[29] = 32'h00000000;
assign filter_banks_17[30] = 32'h00000000;
assign filter_banks_17[31] = 32'h00000000;
assign filter_banks_17[32] = 32'h00000000;
assign filter_banks_17[33] = 32'h00000000;
assign filter_banks_17[34] = 32'h00000000;
assign filter_banks_17[35] = 32'h00000000;
assign filter_banks_17[36] = 32'h00000000;
assign filter_banks_17[37] = 32'h00000000;
assign filter_banks_17[38] = 32'h00000000;
assign filter_banks_17[39] = 32'h00000000;
assign filter_banks_17[40] = 32'h00000000;
assign filter_banks_17[41] = 32'h00000000;
assign filter_banks_17[42] = 32'h00000000;
assign filter_banks_17[43] = 32'h00000000;
assign filter_banks_17[44] = 32'h00000000;
assign filter_banks_17[45] = 32'h00000000;
assign filter_banks_17[46] = 32'h00000000;
assign filter_banks_17[47] = 32'h00000000;
assign filter_banks_17[48] = 32'h00000000;
assign filter_banks_17[49] = 32'h00000000;
assign filter_banks_17[50] = 32'h00000000;
assign filter_banks_17[51] = 32'h00000000;
assign filter_banks_17[52] = 32'h00000000;
assign filter_banks_17[53] = 32'h00000000;
assign filter_banks_17[54] = 32'h00000000;
assign filter_banks_17[55] = 32'h00000000;
assign filter_banks_17[56] = 32'h00000000;
assign filter_banks_17[57] = 32'h00000000;
assign filter_banks_17[58] = 32'h00000000;
assign filter_banks_17[59] = 32'h00000000;
assign filter_banks_17[60] = 32'h00000000;
assign filter_banks_17[61] = 32'h00000000;
assign filter_banks_17[62] = 32'h00000000;
assign filter_banks_17[63] = 32'h00000000;
assign filter_banks_17[64] = 32'h00000000;
assign filter_banks_17[65] = 32'h00000000;
assign filter_banks_17[66] = 32'h00000000;
assign filter_banks_17[67] = 32'h00000000;
assign filter_banks_17[68] = 32'h00000000;
assign filter_banks_17[69] = 32'h00000000;
assign filter_banks_17[70] = 32'h00000000;
assign filter_banks_17[71] = 32'h00000000;
assign filter_banks_17[72] = 32'h00000000;
assign filter_banks_17[73] = 32'h00000000;
assign filter_banks_17[74] = 32'h00000000;
assign filter_banks_17[75] = 32'h00000000;
assign filter_banks_17[76] = 32'h00000000;
assign filter_banks_17[77] = 32'h00000000;
assign filter_banks_17[78] = 32'h3dcccccd;
assign filter_banks_17[79] = 32'h3e4ccccd;
assign filter_banks_17[80] = 32'h3e99999a;
assign filter_banks_17[81] = 32'h3ecccccd;
assign filter_banks_17[82] = 32'h3f000000;
assign filter_banks_17[83] = 32'h3f19999a;
assign filter_banks_17[84] = 32'h3f333333;
assign filter_banks_17[85] = 32'h3f4ccccd;
assign filter_banks_17[86] = 32'h3f666666;
assign filter_banks_17[87] = 32'h3f800000;
assign filter_banks_17[88] = 32'h3f666666;
assign filter_banks_17[89] = 32'h3f4ccccd;
assign filter_banks_17[90] = 32'h3f333333;
assign filter_banks_17[91] = 32'h3f19999a;
assign filter_banks_17[92] = 32'h3f000000;
assign filter_banks_17[93] = 32'h3ecccccd;
assign filter_banks_17[94] = 32'h3e99999a;
assign filter_banks_17[95] = 32'h3e4ccccd;
assign filter_banks_17[96] = 32'h3dcccccd;
assign filter_banks_17[97] = 32'h00000000;
assign filter_banks_17[98] = 32'h00000000;
assign filter_banks_17[99] = 32'h00000000;
assign filter_banks_17[100] = 32'h00000000;
assign filter_banks_17[101] = 32'h00000000;
assign filter_banks_17[102] = 32'h00000000;
assign filter_banks_17[103] = 32'h00000000;
assign filter_banks_17[104] = 32'h00000000;
assign filter_banks_17[105] = 32'h00000000;
assign filter_banks_17[106] = 32'h00000000;
assign filter_banks_17[107] = 32'h00000000;
assign filter_banks_17[108] = 32'h00000000;
assign filter_banks_17[109] = 32'h00000000;
assign filter_banks_17[110] = 32'h00000000;
assign filter_banks_17[111] = 32'h00000000;
assign filter_banks_17[112] = 32'h00000000;
assign filter_banks_17[113] = 32'h00000000;
assign filter_banks_17[114] = 32'h00000000;
assign filter_banks_17[115] = 32'h00000000;
assign filter_banks_17[116] = 32'h00000000;
assign filter_banks_17[117] = 32'h00000000;
assign filter_banks_17[118] = 32'h00000000;
assign filter_banks_17[119] = 32'h00000000;
assign filter_banks_17[120] = 32'h00000000;
assign filter_banks_17[121] = 32'h00000000;
assign filter_banks_17[122] = 32'h00000000;
assign filter_banks_17[123] = 32'h00000000;
assign filter_banks_17[124] = 32'h00000000;
assign filter_banks_17[125] = 32'h00000000;
assign filter_banks_17[126] = 32'h00000000;
assign filter_banks_17[127] = 32'h00000000;
assign filter_banks_17[128] = 32'h00000000;
assign filter_banks_17[129] = 32'h00000000;
assign filter_banks_17[130] = 32'h00000000;
assign filter_banks_17[131] = 32'h00000000;
assign filter_banks_17[132] = 32'h00000000;
assign filter_banks_17[133] = 32'h00000000;
assign filter_banks_17[134] = 32'h00000000;
assign filter_banks_17[135] = 32'h00000000;
assign filter_banks_17[136] = 32'h00000000;
assign filter_banks_17[137] = 32'h00000000;
assign filter_banks_17[138] = 32'h00000000;
assign filter_banks_17[139] = 32'h00000000;
assign filter_banks_17[140] = 32'h00000000;
assign filter_banks_17[141] = 32'h00000000;
assign filter_banks_17[142] = 32'h00000000;
assign filter_banks_17[143] = 32'h00000000;
assign filter_banks_17[144] = 32'h00000000;
assign filter_banks_17[145] = 32'h00000000;
assign filter_banks_17[146] = 32'h00000000;
assign filter_banks_17[147] = 32'h00000000;
assign filter_banks_17[148] = 32'h00000000;
assign filter_banks_17[149] = 32'h00000000;
assign filter_banks_17[150] = 32'h00000000;
assign filter_banks_17[151] = 32'h00000000;
assign filter_banks_17[152] = 32'h00000000;
assign filter_banks_17[153] = 32'h00000000;
assign filter_banks_17[154] = 32'h00000000;
assign filter_banks_17[155] = 32'h00000000;
assign filter_banks_17[156] = 32'h00000000;
assign filter_banks_17[157] = 32'h00000000;
assign filter_banks_17[158] = 32'h00000000;
assign filter_banks_17[159] = 32'h00000000;
assign filter_banks_17[160] = 32'h00000000;
assign filter_banks_17[161] = 32'h00000000;
assign filter_banks_17[162] = 32'h00000000;
assign filter_banks_17[163] = 32'h00000000;
assign filter_banks_17[164] = 32'h00000000;
assign filter_banks_17[165] = 32'h00000000;
assign filter_banks_17[166] = 32'h00000000;
assign filter_banks_17[167] = 32'h00000000;
assign filter_banks_17[168] = 32'h00000000;
assign filter_banks_17[169] = 32'h00000000;
assign filter_banks_17[170] = 32'h00000000;
assign filter_banks_17[171] = 32'h00000000;
assign filter_banks_17[172] = 32'h00000000;
assign filter_banks_17[173] = 32'h00000000;
assign filter_banks_17[174] = 32'h00000000;
assign filter_banks_17[175] = 32'h00000000;
assign filter_banks_17[176] = 32'h00000000;
assign filter_banks_17[177] = 32'h00000000;
assign filter_banks_17[178] = 32'h00000000;
assign filter_banks_17[179] = 32'h00000000;
assign filter_banks_17[180] = 32'h00000000;
assign filter_banks_17[181] = 32'h00000000;
assign filter_banks_17[182] = 32'h00000000;
assign filter_banks_17[183] = 32'h00000000;
assign filter_banks_17[184] = 32'h00000000;
assign filter_banks_17[185] = 32'h00000000;
assign filter_banks_17[186] = 32'h00000000;
assign filter_banks_17[187] = 32'h00000000;
assign filter_banks_17[188] = 32'h00000000;
assign filter_banks_17[189] = 32'h00000000;
assign filter_banks_17[190] = 32'h00000000;
assign filter_banks_17[191] = 32'h00000000;
assign filter_banks_17[192] = 32'h00000000;
assign filter_banks_17[193] = 32'h00000000;
assign filter_banks_17[194] = 32'h00000000;
assign filter_banks_17[195] = 32'h00000000;
assign filter_banks_17[196] = 32'h00000000;
assign filter_banks_17[197] = 32'h00000000;
assign filter_banks_17[198] = 32'h00000000;
assign filter_banks_17[199] = 32'h00000000;
assign filter_banks_17[200] = 32'h00000000;
assign filter_banks_17[201] = 32'h00000000;
assign filter_banks_17[202] = 32'h00000000;
assign filter_banks_17[203] = 32'h00000000;
assign filter_banks_17[204] = 32'h00000000;
assign filter_banks_17[205] = 32'h00000000;
assign filter_banks_17[206] = 32'h00000000;
assign filter_banks_17[207] = 32'h00000000;
assign filter_banks_17[208] = 32'h00000000;
assign filter_banks_17[209] = 32'h00000000;
assign filter_banks_17[210] = 32'h00000000;
assign filter_banks_17[211] = 32'h00000000;
assign filter_banks_17[212] = 32'h00000000;
assign filter_banks_17[213] = 32'h00000000;
assign filter_banks_17[214] = 32'h00000000;
assign filter_banks_17[215] = 32'h00000000;
assign filter_banks_17[216] = 32'h00000000;
assign filter_banks_17[217] = 32'h00000000;
assign filter_banks_17[218] = 32'h00000000;
assign filter_banks_17[219] = 32'h00000000;
assign filter_banks_17[220] = 32'h00000000;
assign filter_banks_17[221] = 32'h00000000;
assign filter_banks_17[222] = 32'h00000000;
assign filter_banks_17[223] = 32'h00000000;
assign filter_banks_17[224] = 32'h00000000;
assign filter_banks_17[225] = 32'h00000000;
assign filter_banks_17[226] = 32'h00000000;
assign filter_banks_17[227] = 32'h00000000;
assign filter_banks_17[228] = 32'h00000000;
assign filter_banks_17[229] = 32'h00000000;
assign filter_banks_17[230] = 32'h00000000;
assign filter_banks_17[231] = 32'h00000000;
assign filter_banks_17[232] = 32'h00000000;
assign filter_banks_17[233] = 32'h00000000;
assign filter_banks_17[234] = 32'h00000000;
assign filter_banks_17[235] = 32'h00000000;
assign filter_banks_17[236] = 32'h00000000;
assign filter_banks_17[237] = 32'h00000000;
assign filter_banks_17[238] = 32'h00000000;
assign filter_banks_17[239] = 32'h00000000;
assign filter_banks_17[240] = 32'h00000000;
assign filter_banks_17[241] = 32'h00000000;
assign filter_banks_17[242] = 32'h00000000;
assign filter_banks_17[243] = 32'h00000000;
assign filter_banks_17[244] = 32'h00000000;
assign filter_banks_17[245] = 32'h00000000;
assign filter_banks_17[246] = 32'h00000000;
assign filter_banks_17[247] = 32'h00000000;
assign filter_banks_17[248] = 32'h00000000;
assign filter_banks_17[249] = 32'h00000000;
assign filter_banks_17[250] = 32'h00000000;
assign filter_banks_17[251] = 32'h00000000;
assign filter_banks_17[252] = 32'h00000000;
assign filter_banks_17[253] = 32'h00000000;
assign filter_banks_17[254] = 32'h00000000;
assign filter_banks_17[255] = 32'h00000000;
assign filter_banks_17[256] = 32'h00000000;
assign filter_banks_18[0] = 32'h00000000;
assign filter_banks_18[1] = 32'h00000000;
assign filter_banks_18[2] = 32'h00000000;
assign filter_banks_18[3] = 32'h00000000;
assign filter_banks_18[4] = 32'h00000000;
assign filter_banks_18[5] = 32'h00000000;
assign filter_banks_18[6] = 32'h00000000;
assign filter_banks_18[7] = 32'h00000000;
assign filter_banks_18[8] = 32'h00000000;
assign filter_banks_18[9] = 32'h00000000;
assign filter_banks_18[10] = 32'h00000000;
assign filter_banks_18[11] = 32'h00000000;
assign filter_banks_18[12] = 32'h00000000;
assign filter_banks_18[13] = 32'h00000000;
assign filter_banks_18[14] = 32'h00000000;
assign filter_banks_18[15] = 32'h00000000;
assign filter_banks_18[16] = 32'h00000000;
assign filter_banks_18[17] = 32'h00000000;
assign filter_banks_18[18] = 32'h00000000;
assign filter_banks_18[19] = 32'h00000000;
assign filter_banks_18[20] = 32'h00000000;
assign filter_banks_18[21] = 32'h00000000;
assign filter_banks_18[22] = 32'h00000000;
assign filter_banks_18[23] = 32'h00000000;
assign filter_banks_18[24] = 32'h00000000;
assign filter_banks_18[25] = 32'h00000000;
assign filter_banks_18[26] = 32'h00000000;
assign filter_banks_18[27] = 32'h00000000;
assign filter_banks_18[28] = 32'h00000000;
assign filter_banks_18[29] = 32'h00000000;
assign filter_banks_18[30] = 32'h00000000;
assign filter_banks_18[31] = 32'h00000000;
assign filter_banks_18[32] = 32'h00000000;
assign filter_banks_18[33] = 32'h00000000;
assign filter_banks_18[34] = 32'h00000000;
assign filter_banks_18[35] = 32'h00000000;
assign filter_banks_18[36] = 32'h00000000;
assign filter_banks_18[37] = 32'h00000000;
assign filter_banks_18[38] = 32'h00000000;
assign filter_banks_18[39] = 32'h00000000;
assign filter_banks_18[40] = 32'h00000000;
assign filter_banks_18[41] = 32'h00000000;
assign filter_banks_18[42] = 32'h00000000;
assign filter_banks_18[43] = 32'h00000000;
assign filter_banks_18[44] = 32'h00000000;
assign filter_banks_18[45] = 32'h00000000;
assign filter_banks_18[46] = 32'h00000000;
assign filter_banks_18[47] = 32'h00000000;
assign filter_banks_18[48] = 32'h00000000;
assign filter_banks_18[49] = 32'h00000000;
assign filter_banks_18[50] = 32'h00000000;
assign filter_banks_18[51] = 32'h00000000;
assign filter_banks_18[52] = 32'h00000000;
assign filter_banks_18[53] = 32'h00000000;
assign filter_banks_18[54] = 32'h00000000;
assign filter_banks_18[55] = 32'h00000000;
assign filter_banks_18[56] = 32'h00000000;
assign filter_banks_18[57] = 32'h00000000;
assign filter_banks_18[58] = 32'h00000000;
assign filter_banks_18[59] = 32'h00000000;
assign filter_banks_18[60] = 32'h00000000;
assign filter_banks_18[61] = 32'h00000000;
assign filter_banks_18[62] = 32'h00000000;
assign filter_banks_18[63] = 32'h00000000;
assign filter_banks_18[64] = 32'h00000000;
assign filter_banks_18[65] = 32'h00000000;
assign filter_banks_18[66] = 32'h00000000;
assign filter_banks_18[67] = 32'h00000000;
assign filter_banks_18[68] = 32'h00000000;
assign filter_banks_18[69] = 32'h00000000;
assign filter_banks_18[70] = 32'h00000000;
assign filter_banks_18[71] = 32'h00000000;
assign filter_banks_18[72] = 32'h00000000;
assign filter_banks_18[73] = 32'h00000000;
assign filter_banks_18[74] = 32'h00000000;
assign filter_banks_18[75] = 32'h00000000;
assign filter_banks_18[76] = 32'h00000000;
assign filter_banks_18[77] = 32'h00000000;
assign filter_banks_18[78] = 32'h00000000;
assign filter_banks_18[79] = 32'h00000000;
assign filter_banks_18[80] = 32'h00000000;
assign filter_banks_18[81] = 32'h00000000;
assign filter_banks_18[82] = 32'h00000000;
assign filter_banks_18[83] = 32'h00000000;
assign filter_banks_18[84] = 32'h00000000;
assign filter_banks_18[85] = 32'h00000000;
assign filter_banks_18[86] = 32'h00000000;
assign filter_banks_18[87] = 32'h00000000;
assign filter_banks_18[88] = 32'h3dcccccd;
assign filter_banks_18[89] = 32'h3e4ccccd;
assign filter_banks_18[90] = 32'h3e99999a;
assign filter_banks_18[91] = 32'h3ecccccd;
assign filter_banks_18[92] = 32'h3f000000;
assign filter_banks_18[93] = 32'h3f19999a;
assign filter_banks_18[94] = 32'h3f333333;
assign filter_banks_18[95] = 32'h3f4ccccd;
assign filter_banks_18[96] = 32'h3f666666;
assign filter_banks_18[97] = 32'h3f800000;
assign filter_banks_18[98] = 32'h3f6aaaab;
assign filter_banks_18[99] = 32'h3f555555;
assign filter_banks_18[100] = 32'h3f400000;
assign filter_banks_18[101] = 32'h3f2aaaab;
assign filter_banks_18[102] = 32'h3f155555;
assign filter_banks_18[103] = 32'h3f000000;
assign filter_banks_18[104] = 32'h3ed55555;
assign filter_banks_18[105] = 32'h3eaaaaab;
assign filter_banks_18[106] = 32'h3e800000;
assign filter_banks_18[107] = 32'h3e2aaaab;
assign filter_banks_18[108] = 32'h3daaaaab;
assign filter_banks_18[109] = 32'h00000000;
assign filter_banks_18[110] = 32'h00000000;
assign filter_banks_18[111] = 32'h00000000;
assign filter_banks_18[112] = 32'h00000000;
assign filter_banks_18[113] = 32'h00000000;
assign filter_banks_18[114] = 32'h00000000;
assign filter_banks_18[115] = 32'h00000000;
assign filter_banks_18[116] = 32'h00000000;
assign filter_banks_18[117] = 32'h00000000;
assign filter_banks_18[118] = 32'h00000000;
assign filter_banks_18[119] = 32'h00000000;
assign filter_banks_18[120] = 32'h00000000;
assign filter_banks_18[121] = 32'h00000000;
assign filter_banks_18[122] = 32'h00000000;
assign filter_banks_18[123] = 32'h00000000;
assign filter_banks_18[124] = 32'h00000000;
assign filter_banks_18[125] = 32'h00000000;
assign filter_banks_18[126] = 32'h00000000;
assign filter_banks_18[127] = 32'h00000000;
assign filter_banks_18[128] = 32'h00000000;
assign filter_banks_18[129] = 32'h00000000;
assign filter_banks_18[130] = 32'h00000000;
assign filter_banks_18[131] = 32'h00000000;
assign filter_banks_18[132] = 32'h00000000;
assign filter_banks_18[133] = 32'h00000000;
assign filter_banks_18[134] = 32'h00000000;
assign filter_banks_18[135] = 32'h00000000;
assign filter_banks_18[136] = 32'h00000000;
assign filter_banks_18[137] = 32'h00000000;
assign filter_banks_18[138] = 32'h00000000;
assign filter_banks_18[139] = 32'h00000000;
assign filter_banks_18[140] = 32'h00000000;
assign filter_banks_18[141] = 32'h00000000;
assign filter_banks_18[142] = 32'h00000000;
assign filter_banks_18[143] = 32'h00000000;
assign filter_banks_18[144] = 32'h00000000;
assign filter_banks_18[145] = 32'h00000000;
assign filter_banks_18[146] = 32'h00000000;
assign filter_banks_18[147] = 32'h00000000;
assign filter_banks_18[148] = 32'h00000000;
assign filter_banks_18[149] = 32'h00000000;
assign filter_banks_18[150] = 32'h00000000;
assign filter_banks_18[151] = 32'h00000000;
assign filter_banks_18[152] = 32'h00000000;
assign filter_banks_18[153] = 32'h00000000;
assign filter_banks_18[154] = 32'h00000000;
assign filter_banks_18[155] = 32'h00000000;
assign filter_banks_18[156] = 32'h00000000;
assign filter_banks_18[157] = 32'h00000000;
assign filter_banks_18[158] = 32'h00000000;
assign filter_banks_18[159] = 32'h00000000;
assign filter_banks_18[160] = 32'h00000000;
assign filter_banks_18[161] = 32'h00000000;
assign filter_banks_18[162] = 32'h00000000;
assign filter_banks_18[163] = 32'h00000000;
assign filter_banks_18[164] = 32'h00000000;
assign filter_banks_18[165] = 32'h00000000;
assign filter_banks_18[166] = 32'h00000000;
assign filter_banks_18[167] = 32'h00000000;
assign filter_banks_18[168] = 32'h00000000;
assign filter_banks_18[169] = 32'h00000000;
assign filter_banks_18[170] = 32'h00000000;
assign filter_banks_18[171] = 32'h00000000;
assign filter_banks_18[172] = 32'h00000000;
assign filter_banks_18[173] = 32'h00000000;
assign filter_banks_18[174] = 32'h00000000;
assign filter_banks_18[175] = 32'h00000000;
assign filter_banks_18[176] = 32'h00000000;
assign filter_banks_18[177] = 32'h00000000;
assign filter_banks_18[178] = 32'h00000000;
assign filter_banks_18[179] = 32'h00000000;
assign filter_banks_18[180] = 32'h00000000;
assign filter_banks_18[181] = 32'h00000000;
assign filter_banks_18[182] = 32'h00000000;
assign filter_banks_18[183] = 32'h00000000;
assign filter_banks_18[184] = 32'h00000000;
assign filter_banks_18[185] = 32'h00000000;
assign filter_banks_18[186] = 32'h00000000;
assign filter_banks_18[187] = 32'h00000000;
assign filter_banks_18[188] = 32'h00000000;
assign filter_banks_18[189] = 32'h00000000;
assign filter_banks_18[190] = 32'h00000000;
assign filter_banks_18[191] = 32'h00000000;
assign filter_banks_18[192] = 32'h00000000;
assign filter_banks_18[193] = 32'h00000000;
assign filter_banks_18[194] = 32'h00000000;
assign filter_banks_18[195] = 32'h00000000;
assign filter_banks_18[196] = 32'h00000000;
assign filter_banks_18[197] = 32'h00000000;
assign filter_banks_18[198] = 32'h00000000;
assign filter_banks_18[199] = 32'h00000000;
assign filter_banks_18[200] = 32'h00000000;
assign filter_banks_18[201] = 32'h00000000;
assign filter_banks_18[202] = 32'h00000000;
assign filter_banks_18[203] = 32'h00000000;
assign filter_banks_18[204] = 32'h00000000;
assign filter_banks_18[205] = 32'h00000000;
assign filter_banks_18[206] = 32'h00000000;
assign filter_banks_18[207] = 32'h00000000;
assign filter_banks_18[208] = 32'h00000000;
assign filter_banks_18[209] = 32'h00000000;
assign filter_banks_18[210] = 32'h00000000;
assign filter_banks_18[211] = 32'h00000000;
assign filter_banks_18[212] = 32'h00000000;
assign filter_banks_18[213] = 32'h00000000;
assign filter_banks_18[214] = 32'h00000000;
assign filter_banks_18[215] = 32'h00000000;
assign filter_banks_18[216] = 32'h00000000;
assign filter_banks_18[217] = 32'h00000000;
assign filter_banks_18[218] = 32'h00000000;
assign filter_banks_18[219] = 32'h00000000;
assign filter_banks_18[220] = 32'h00000000;
assign filter_banks_18[221] = 32'h00000000;
assign filter_banks_18[222] = 32'h00000000;
assign filter_banks_18[223] = 32'h00000000;
assign filter_banks_18[224] = 32'h00000000;
assign filter_banks_18[225] = 32'h00000000;
assign filter_banks_18[226] = 32'h00000000;
assign filter_banks_18[227] = 32'h00000000;
assign filter_banks_18[228] = 32'h00000000;
assign filter_banks_18[229] = 32'h00000000;
assign filter_banks_18[230] = 32'h00000000;
assign filter_banks_18[231] = 32'h00000000;
assign filter_banks_18[232] = 32'h00000000;
assign filter_banks_18[233] = 32'h00000000;
assign filter_banks_18[234] = 32'h00000000;
assign filter_banks_18[235] = 32'h00000000;
assign filter_banks_18[236] = 32'h00000000;
assign filter_banks_18[237] = 32'h00000000;
assign filter_banks_18[238] = 32'h00000000;
assign filter_banks_18[239] = 32'h00000000;
assign filter_banks_18[240] = 32'h00000000;
assign filter_banks_18[241] = 32'h00000000;
assign filter_banks_18[242] = 32'h00000000;
assign filter_banks_18[243] = 32'h00000000;
assign filter_banks_18[244] = 32'h00000000;
assign filter_banks_18[245] = 32'h00000000;
assign filter_banks_18[246] = 32'h00000000;
assign filter_banks_18[247] = 32'h00000000;
assign filter_banks_18[248] = 32'h00000000;
assign filter_banks_18[249] = 32'h00000000;
assign filter_banks_18[250] = 32'h00000000;
assign filter_banks_18[251] = 32'h00000000;
assign filter_banks_18[252] = 32'h00000000;
assign filter_banks_18[253] = 32'h00000000;
assign filter_banks_18[254] = 32'h00000000;
assign filter_banks_18[255] = 32'h00000000;
assign filter_banks_18[256] = 32'h00000000;
assign filter_banks_19[0] = 32'h00000000;
assign filter_banks_19[1] = 32'h00000000;
assign filter_banks_19[2] = 32'h00000000;
assign filter_banks_19[3] = 32'h00000000;
assign filter_banks_19[4] = 32'h00000000;
assign filter_banks_19[5] = 32'h00000000;
assign filter_banks_19[6] = 32'h00000000;
assign filter_banks_19[7] = 32'h00000000;
assign filter_banks_19[8] = 32'h00000000;
assign filter_banks_19[9] = 32'h00000000;
assign filter_banks_19[10] = 32'h00000000;
assign filter_banks_19[11] = 32'h00000000;
assign filter_banks_19[12] = 32'h00000000;
assign filter_banks_19[13] = 32'h00000000;
assign filter_banks_19[14] = 32'h00000000;
assign filter_banks_19[15] = 32'h00000000;
assign filter_banks_19[16] = 32'h00000000;
assign filter_banks_19[17] = 32'h00000000;
assign filter_banks_19[18] = 32'h00000000;
assign filter_banks_19[19] = 32'h00000000;
assign filter_banks_19[20] = 32'h00000000;
assign filter_banks_19[21] = 32'h00000000;
assign filter_banks_19[22] = 32'h00000000;
assign filter_banks_19[23] = 32'h00000000;
assign filter_banks_19[24] = 32'h00000000;
assign filter_banks_19[25] = 32'h00000000;
assign filter_banks_19[26] = 32'h00000000;
assign filter_banks_19[27] = 32'h00000000;
assign filter_banks_19[28] = 32'h00000000;
assign filter_banks_19[29] = 32'h00000000;
assign filter_banks_19[30] = 32'h00000000;
assign filter_banks_19[31] = 32'h00000000;
assign filter_banks_19[32] = 32'h00000000;
assign filter_banks_19[33] = 32'h00000000;
assign filter_banks_19[34] = 32'h00000000;
assign filter_banks_19[35] = 32'h00000000;
assign filter_banks_19[36] = 32'h00000000;
assign filter_banks_19[37] = 32'h00000000;
assign filter_banks_19[38] = 32'h00000000;
assign filter_banks_19[39] = 32'h00000000;
assign filter_banks_19[40] = 32'h00000000;
assign filter_banks_19[41] = 32'h00000000;
assign filter_banks_19[42] = 32'h00000000;
assign filter_banks_19[43] = 32'h00000000;
assign filter_banks_19[44] = 32'h00000000;
assign filter_banks_19[45] = 32'h00000000;
assign filter_banks_19[46] = 32'h00000000;
assign filter_banks_19[47] = 32'h00000000;
assign filter_banks_19[48] = 32'h00000000;
assign filter_banks_19[49] = 32'h00000000;
assign filter_banks_19[50] = 32'h00000000;
assign filter_banks_19[51] = 32'h00000000;
assign filter_banks_19[52] = 32'h00000000;
assign filter_banks_19[53] = 32'h00000000;
assign filter_banks_19[54] = 32'h00000000;
assign filter_banks_19[55] = 32'h00000000;
assign filter_banks_19[56] = 32'h00000000;
assign filter_banks_19[57] = 32'h00000000;
assign filter_banks_19[58] = 32'h00000000;
assign filter_banks_19[59] = 32'h00000000;
assign filter_banks_19[60] = 32'h00000000;
assign filter_banks_19[61] = 32'h00000000;
assign filter_banks_19[62] = 32'h00000000;
assign filter_banks_19[63] = 32'h00000000;
assign filter_banks_19[64] = 32'h00000000;
assign filter_banks_19[65] = 32'h00000000;
assign filter_banks_19[66] = 32'h00000000;
assign filter_banks_19[67] = 32'h00000000;
assign filter_banks_19[68] = 32'h00000000;
assign filter_banks_19[69] = 32'h00000000;
assign filter_banks_19[70] = 32'h00000000;
assign filter_banks_19[71] = 32'h00000000;
assign filter_banks_19[72] = 32'h00000000;
assign filter_banks_19[73] = 32'h00000000;
assign filter_banks_19[74] = 32'h00000000;
assign filter_banks_19[75] = 32'h00000000;
assign filter_banks_19[76] = 32'h00000000;
assign filter_banks_19[77] = 32'h00000000;
assign filter_banks_19[78] = 32'h00000000;
assign filter_banks_19[79] = 32'h00000000;
assign filter_banks_19[80] = 32'h00000000;
assign filter_banks_19[81] = 32'h00000000;
assign filter_banks_19[82] = 32'h00000000;
assign filter_banks_19[83] = 32'h00000000;
assign filter_banks_19[84] = 32'h00000000;
assign filter_banks_19[85] = 32'h00000000;
assign filter_banks_19[86] = 32'h00000000;
assign filter_banks_19[87] = 32'h00000000;
assign filter_banks_19[88] = 32'h00000000;
assign filter_banks_19[89] = 32'h00000000;
assign filter_banks_19[90] = 32'h00000000;
assign filter_banks_19[91] = 32'h00000000;
assign filter_banks_19[92] = 32'h00000000;
assign filter_banks_19[93] = 32'h00000000;
assign filter_banks_19[94] = 32'h00000000;
assign filter_banks_19[95] = 32'h00000000;
assign filter_banks_19[96] = 32'h00000000;
assign filter_banks_19[97] = 32'h00000000;
assign filter_banks_19[98] = 32'h3daaaaab;
assign filter_banks_19[99] = 32'h3e2aaaab;
assign filter_banks_19[100] = 32'h3e800000;
assign filter_banks_19[101] = 32'h3eaaaaab;
assign filter_banks_19[102] = 32'h3ed55555;
assign filter_banks_19[103] = 32'h3f000000;
assign filter_banks_19[104] = 32'h3f155555;
assign filter_banks_19[105] = 32'h3f2aaaab;
assign filter_banks_19[106] = 32'h3f400000;
assign filter_banks_19[107] = 32'h3f555555;
assign filter_banks_19[108] = 32'h3f6aaaab;
assign filter_banks_19[109] = 32'h3f800000;
assign filter_banks_19[110] = 32'h3f6c4ec5;
assign filter_banks_19[111] = 32'h3f589d8a;
assign filter_banks_19[112] = 32'h3f44ec4f;
assign filter_banks_19[113] = 32'h3f313b14;
assign filter_banks_19[114] = 32'h3f1d89d9;
assign filter_banks_19[115] = 32'h3f09d89e;
assign filter_banks_19[116] = 32'h3eec4ec5;
assign filter_banks_19[117] = 32'h3ec4ec4f;
assign filter_banks_19[118] = 32'h3e9d89d9;
assign filter_banks_19[119] = 32'h3e6c4ec5;
assign filter_banks_19[120] = 32'h3e1d89d9;
assign filter_banks_19[121] = 32'h3d9d89d9;
assign filter_banks_19[122] = 32'h00000000;
assign filter_banks_19[123] = 32'h00000000;
assign filter_banks_19[124] = 32'h00000000;
assign filter_banks_19[125] = 32'h00000000;
assign filter_banks_19[126] = 32'h00000000;
assign filter_banks_19[127] = 32'h00000000;
assign filter_banks_19[128] = 32'h00000000;
assign filter_banks_19[129] = 32'h00000000;
assign filter_banks_19[130] = 32'h00000000;
assign filter_banks_19[131] = 32'h00000000;
assign filter_banks_19[132] = 32'h00000000;
assign filter_banks_19[133] = 32'h00000000;
assign filter_banks_19[134] = 32'h00000000;
assign filter_banks_19[135] = 32'h00000000;
assign filter_banks_19[136] = 32'h00000000;
assign filter_banks_19[137] = 32'h00000000;
assign filter_banks_19[138] = 32'h00000000;
assign filter_banks_19[139] = 32'h00000000;
assign filter_banks_19[140] = 32'h00000000;
assign filter_banks_19[141] = 32'h00000000;
assign filter_banks_19[142] = 32'h00000000;
assign filter_banks_19[143] = 32'h00000000;
assign filter_banks_19[144] = 32'h00000000;
assign filter_banks_19[145] = 32'h00000000;
assign filter_banks_19[146] = 32'h00000000;
assign filter_banks_19[147] = 32'h00000000;
assign filter_banks_19[148] = 32'h00000000;
assign filter_banks_19[149] = 32'h00000000;
assign filter_banks_19[150] = 32'h00000000;
assign filter_banks_19[151] = 32'h00000000;
assign filter_banks_19[152] = 32'h00000000;
assign filter_banks_19[153] = 32'h00000000;
assign filter_banks_19[154] = 32'h00000000;
assign filter_banks_19[155] = 32'h00000000;
assign filter_banks_19[156] = 32'h00000000;
assign filter_banks_19[157] = 32'h00000000;
assign filter_banks_19[158] = 32'h00000000;
assign filter_banks_19[159] = 32'h00000000;
assign filter_banks_19[160] = 32'h00000000;
assign filter_banks_19[161] = 32'h00000000;
assign filter_banks_19[162] = 32'h00000000;
assign filter_banks_19[163] = 32'h00000000;
assign filter_banks_19[164] = 32'h00000000;
assign filter_banks_19[165] = 32'h00000000;
assign filter_banks_19[166] = 32'h00000000;
assign filter_banks_19[167] = 32'h00000000;
assign filter_banks_19[168] = 32'h00000000;
assign filter_banks_19[169] = 32'h00000000;
assign filter_banks_19[170] = 32'h00000000;
assign filter_banks_19[171] = 32'h00000000;
assign filter_banks_19[172] = 32'h00000000;
assign filter_banks_19[173] = 32'h00000000;
assign filter_banks_19[174] = 32'h00000000;
assign filter_banks_19[175] = 32'h00000000;
assign filter_banks_19[176] = 32'h00000000;
assign filter_banks_19[177] = 32'h00000000;
assign filter_banks_19[178] = 32'h00000000;
assign filter_banks_19[179] = 32'h00000000;
assign filter_banks_19[180] = 32'h00000000;
assign filter_banks_19[181] = 32'h00000000;
assign filter_banks_19[182] = 32'h00000000;
assign filter_banks_19[183] = 32'h00000000;
assign filter_banks_19[184] = 32'h00000000;
assign filter_banks_19[185] = 32'h00000000;
assign filter_banks_19[186] = 32'h00000000;
assign filter_banks_19[187] = 32'h00000000;
assign filter_banks_19[188] = 32'h00000000;
assign filter_banks_19[189] = 32'h00000000;
assign filter_banks_19[190] = 32'h00000000;
assign filter_banks_19[191] = 32'h00000000;
assign filter_banks_19[192] = 32'h00000000;
assign filter_banks_19[193] = 32'h00000000;
assign filter_banks_19[194] = 32'h00000000;
assign filter_banks_19[195] = 32'h00000000;
assign filter_banks_19[196] = 32'h00000000;
assign filter_banks_19[197] = 32'h00000000;
assign filter_banks_19[198] = 32'h00000000;
assign filter_banks_19[199] = 32'h00000000;
assign filter_banks_19[200] = 32'h00000000;
assign filter_banks_19[201] = 32'h00000000;
assign filter_banks_19[202] = 32'h00000000;
assign filter_banks_19[203] = 32'h00000000;
assign filter_banks_19[204] = 32'h00000000;
assign filter_banks_19[205] = 32'h00000000;
assign filter_banks_19[206] = 32'h00000000;
assign filter_banks_19[207] = 32'h00000000;
assign filter_banks_19[208] = 32'h00000000;
assign filter_banks_19[209] = 32'h00000000;
assign filter_banks_19[210] = 32'h00000000;
assign filter_banks_19[211] = 32'h00000000;
assign filter_banks_19[212] = 32'h00000000;
assign filter_banks_19[213] = 32'h00000000;
assign filter_banks_19[214] = 32'h00000000;
assign filter_banks_19[215] = 32'h00000000;
assign filter_banks_19[216] = 32'h00000000;
assign filter_banks_19[217] = 32'h00000000;
assign filter_banks_19[218] = 32'h00000000;
assign filter_banks_19[219] = 32'h00000000;
assign filter_banks_19[220] = 32'h00000000;
assign filter_banks_19[221] = 32'h00000000;
assign filter_banks_19[222] = 32'h00000000;
assign filter_banks_19[223] = 32'h00000000;
assign filter_banks_19[224] = 32'h00000000;
assign filter_banks_19[225] = 32'h00000000;
assign filter_banks_19[226] = 32'h00000000;
assign filter_banks_19[227] = 32'h00000000;
assign filter_banks_19[228] = 32'h00000000;
assign filter_banks_19[229] = 32'h00000000;
assign filter_banks_19[230] = 32'h00000000;
assign filter_banks_19[231] = 32'h00000000;
assign filter_banks_19[232] = 32'h00000000;
assign filter_banks_19[233] = 32'h00000000;
assign filter_banks_19[234] = 32'h00000000;
assign filter_banks_19[235] = 32'h00000000;
assign filter_banks_19[236] = 32'h00000000;
assign filter_banks_19[237] = 32'h00000000;
assign filter_banks_19[238] = 32'h00000000;
assign filter_banks_19[239] = 32'h00000000;
assign filter_banks_19[240] = 32'h00000000;
assign filter_banks_19[241] = 32'h00000000;
assign filter_banks_19[242] = 32'h00000000;
assign filter_banks_19[243] = 32'h00000000;
assign filter_banks_19[244] = 32'h00000000;
assign filter_banks_19[245] = 32'h00000000;
assign filter_banks_19[246] = 32'h00000000;
assign filter_banks_19[247] = 32'h00000000;
assign filter_banks_19[248] = 32'h00000000;
assign filter_banks_19[249] = 32'h00000000;
assign filter_banks_19[250] = 32'h00000000;
assign filter_banks_19[251] = 32'h00000000;
assign filter_banks_19[252] = 32'h00000000;
assign filter_banks_19[253] = 32'h00000000;
assign filter_banks_19[254] = 32'h00000000;
assign filter_banks_19[255] = 32'h00000000;
assign filter_banks_19[256] = 32'h00000000;
assign filter_banks_20[0] = 32'h00000000;
assign filter_banks_20[1] = 32'h00000000;
assign filter_banks_20[2] = 32'h00000000;
assign filter_banks_20[3] = 32'h00000000;
assign filter_banks_20[4] = 32'h00000000;
assign filter_banks_20[5] = 32'h00000000;
assign filter_banks_20[6] = 32'h00000000;
assign filter_banks_20[7] = 32'h00000000;
assign filter_banks_20[8] = 32'h00000000;
assign filter_banks_20[9] = 32'h00000000;
assign filter_banks_20[10] = 32'h00000000;
assign filter_banks_20[11] = 32'h00000000;
assign filter_banks_20[12] = 32'h00000000;
assign filter_banks_20[13] = 32'h00000000;
assign filter_banks_20[14] = 32'h00000000;
assign filter_banks_20[15] = 32'h00000000;
assign filter_banks_20[16] = 32'h00000000;
assign filter_banks_20[17] = 32'h00000000;
assign filter_banks_20[18] = 32'h00000000;
assign filter_banks_20[19] = 32'h00000000;
assign filter_banks_20[20] = 32'h00000000;
assign filter_banks_20[21] = 32'h00000000;
assign filter_banks_20[22] = 32'h00000000;
assign filter_banks_20[23] = 32'h00000000;
assign filter_banks_20[24] = 32'h00000000;
assign filter_banks_20[25] = 32'h00000000;
assign filter_banks_20[26] = 32'h00000000;
assign filter_banks_20[27] = 32'h00000000;
assign filter_banks_20[28] = 32'h00000000;
assign filter_banks_20[29] = 32'h00000000;
assign filter_banks_20[30] = 32'h00000000;
assign filter_banks_20[31] = 32'h00000000;
assign filter_banks_20[32] = 32'h00000000;
assign filter_banks_20[33] = 32'h00000000;
assign filter_banks_20[34] = 32'h00000000;
assign filter_banks_20[35] = 32'h00000000;
assign filter_banks_20[36] = 32'h00000000;
assign filter_banks_20[37] = 32'h00000000;
assign filter_banks_20[38] = 32'h00000000;
assign filter_banks_20[39] = 32'h00000000;
assign filter_banks_20[40] = 32'h00000000;
assign filter_banks_20[41] = 32'h00000000;
assign filter_banks_20[42] = 32'h00000000;
assign filter_banks_20[43] = 32'h00000000;
assign filter_banks_20[44] = 32'h00000000;
assign filter_banks_20[45] = 32'h00000000;
assign filter_banks_20[46] = 32'h00000000;
assign filter_banks_20[47] = 32'h00000000;
assign filter_banks_20[48] = 32'h00000000;
assign filter_banks_20[49] = 32'h00000000;
assign filter_banks_20[50] = 32'h00000000;
assign filter_banks_20[51] = 32'h00000000;
assign filter_banks_20[52] = 32'h00000000;
assign filter_banks_20[53] = 32'h00000000;
assign filter_banks_20[54] = 32'h00000000;
assign filter_banks_20[55] = 32'h00000000;
assign filter_banks_20[56] = 32'h00000000;
assign filter_banks_20[57] = 32'h00000000;
assign filter_banks_20[58] = 32'h00000000;
assign filter_banks_20[59] = 32'h00000000;
assign filter_banks_20[60] = 32'h00000000;
assign filter_banks_20[61] = 32'h00000000;
assign filter_banks_20[62] = 32'h00000000;
assign filter_banks_20[63] = 32'h00000000;
assign filter_banks_20[64] = 32'h00000000;
assign filter_banks_20[65] = 32'h00000000;
assign filter_banks_20[66] = 32'h00000000;
assign filter_banks_20[67] = 32'h00000000;
assign filter_banks_20[68] = 32'h00000000;
assign filter_banks_20[69] = 32'h00000000;
assign filter_banks_20[70] = 32'h00000000;
assign filter_banks_20[71] = 32'h00000000;
assign filter_banks_20[72] = 32'h00000000;
assign filter_banks_20[73] = 32'h00000000;
assign filter_banks_20[74] = 32'h00000000;
assign filter_banks_20[75] = 32'h00000000;
assign filter_banks_20[76] = 32'h00000000;
assign filter_banks_20[77] = 32'h00000000;
assign filter_banks_20[78] = 32'h00000000;
assign filter_banks_20[79] = 32'h00000000;
assign filter_banks_20[80] = 32'h00000000;
assign filter_banks_20[81] = 32'h00000000;
assign filter_banks_20[82] = 32'h00000000;
assign filter_banks_20[83] = 32'h00000000;
assign filter_banks_20[84] = 32'h00000000;
assign filter_banks_20[85] = 32'h00000000;
assign filter_banks_20[86] = 32'h00000000;
assign filter_banks_20[87] = 32'h00000000;
assign filter_banks_20[88] = 32'h00000000;
assign filter_banks_20[89] = 32'h00000000;
assign filter_banks_20[90] = 32'h00000000;
assign filter_banks_20[91] = 32'h00000000;
assign filter_banks_20[92] = 32'h00000000;
assign filter_banks_20[93] = 32'h00000000;
assign filter_banks_20[94] = 32'h00000000;
assign filter_banks_20[95] = 32'h00000000;
assign filter_banks_20[96] = 32'h00000000;
assign filter_banks_20[97] = 32'h00000000;
assign filter_banks_20[98] = 32'h00000000;
assign filter_banks_20[99] = 32'h00000000;
assign filter_banks_20[100] = 32'h00000000;
assign filter_banks_20[101] = 32'h00000000;
assign filter_banks_20[102] = 32'h00000000;
assign filter_banks_20[103] = 32'h00000000;
assign filter_banks_20[104] = 32'h00000000;
assign filter_banks_20[105] = 32'h00000000;
assign filter_banks_20[106] = 32'h00000000;
assign filter_banks_20[107] = 32'h00000000;
assign filter_banks_20[108] = 32'h00000000;
assign filter_banks_20[109] = 32'h00000000;
assign filter_banks_20[110] = 32'h3d9d89d9;
assign filter_banks_20[111] = 32'h3e1d89d9;
assign filter_banks_20[112] = 32'h3e6c4ec5;
assign filter_banks_20[113] = 32'h3e9d89d9;
assign filter_banks_20[114] = 32'h3ec4ec4f;
assign filter_banks_20[115] = 32'h3eec4ec5;
assign filter_banks_20[116] = 32'h3f09d89e;
assign filter_banks_20[117] = 32'h3f1d89d9;
assign filter_banks_20[118] = 32'h3f313b14;
assign filter_banks_20[119] = 32'h3f44ec4f;
assign filter_banks_20[120] = 32'h3f589d8a;
assign filter_banks_20[121] = 32'h3f6c4ec5;
assign filter_banks_20[122] = 32'h3f800000;
assign filter_banks_20[123] = 32'h3f6db6db;
assign filter_banks_20[124] = 32'h3f5b6db7;
assign filter_banks_20[125] = 32'h3f492492;
assign filter_banks_20[126] = 32'h3f36db6e;
assign filter_banks_20[127] = 32'h3f249249;
assign filter_banks_20[128] = 32'h3f124925;
assign filter_banks_20[129] = 32'h3f000000;
assign filter_banks_20[130] = 32'h3edb6db7;
assign filter_banks_20[131] = 32'h3eb6db6e;
assign filter_banks_20[132] = 32'h3e924925;
assign filter_banks_20[133] = 32'h3e5b6db7;
assign filter_banks_20[134] = 32'h3e124925;
assign filter_banks_20[135] = 32'h3d924925;
assign filter_banks_20[136] = 32'h00000000;
assign filter_banks_20[137] = 32'h00000000;
assign filter_banks_20[138] = 32'h00000000;
assign filter_banks_20[139] = 32'h00000000;
assign filter_banks_20[140] = 32'h00000000;
assign filter_banks_20[141] = 32'h00000000;
assign filter_banks_20[142] = 32'h00000000;
assign filter_banks_20[143] = 32'h00000000;
assign filter_banks_20[144] = 32'h00000000;
assign filter_banks_20[145] = 32'h00000000;
assign filter_banks_20[146] = 32'h00000000;
assign filter_banks_20[147] = 32'h00000000;
assign filter_banks_20[148] = 32'h00000000;
assign filter_banks_20[149] = 32'h00000000;
assign filter_banks_20[150] = 32'h00000000;
assign filter_banks_20[151] = 32'h00000000;
assign filter_banks_20[152] = 32'h00000000;
assign filter_banks_20[153] = 32'h00000000;
assign filter_banks_20[154] = 32'h00000000;
assign filter_banks_20[155] = 32'h00000000;
assign filter_banks_20[156] = 32'h00000000;
assign filter_banks_20[157] = 32'h00000000;
assign filter_banks_20[158] = 32'h00000000;
assign filter_banks_20[159] = 32'h00000000;
assign filter_banks_20[160] = 32'h00000000;
assign filter_banks_20[161] = 32'h00000000;
assign filter_banks_20[162] = 32'h00000000;
assign filter_banks_20[163] = 32'h00000000;
assign filter_banks_20[164] = 32'h00000000;
assign filter_banks_20[165] = 32'h00000000;
assign filter_banks_20[166] = 32'h00000000;
assign filter_banks_20[167] = 32'h00000000;
assign filter_banks_20[168] = 32'h00000000;
assign filter_banks_20[169] = 32'h00000000;
assign filter_banks_20[170] = 32'h00000000;
assign filter_banks_20[171] = 32'h00000000;
assign filter_banks_20[172] = 32'h00000000;
assign filter_banks_20[173] = 32'h00000000;
assign filter_banks_20[174] = 32'h00000000;
assign filter_banks_20[175] = 32'h00000000;
assign filter_banks_20[176] = 32'h00000000;
assign filter_banks_20[177] = 32'h00000000;
assign filter_banks_20[178] = 32'h00000000;
assign filter_banks_20[179] = 32'h00000000;
assign filter_banks_20[180] = 32'h00000000;
assign filter_banks_20[181] = 32'h00000000;
assign filter_banks_20[182] = 32'h00000000;
assign filter_banks_20[183] = 32'h00000000;
assign filter_banks_20[184] = 32'h00000000;
assign filter_banks_20[185] = 32'h00000000;
assign filter_banks_20[186] = 32'h00000000;
assign filter_banks_20[187] = 32'h00000000;
assign filter_banks_20[188] = 32'h00000000;
assign filter_banks_20[189] = 32'h00000000;
assign filter_banks_20[190] = 32'h00000000;
assign filter_banks_20[191] = 32'h00000000;
assign filter_banks_20[192] = 32'h00000000;
assign filter_banks_20[193] = 32'h00000000;
assign filter_banks_20[194] = 32'h00000000;
assign filter_banks_20[195] = 32'h00000000;
assign filter_banks_20[196] = 32'h00000000;
assign filter_banks_20[197] = 32'h00000000;
assign filter_banks_20[198] = 32'h00000000;
assign filter_banks_20[199] = 32'h00000000;
assign filter_banks_20[200] = 32'h00000000;
assign filter_banks_20[201] = 32'h00000000;
assign filter_banks_20[202] = 32'h00000000;
assign filter_banks_20[203] = 32'h00000000;
assign filter_banks_20[204] = 32'h00000000;
assign filter_banks_20[205] = 32'h00000000;
assign filter_banks_20[206] = 32'h00000000;
assign filter_banks_20[207] = 32'h00000000;
assign filter_banks_20[208] = 32'h00000000;
assign filter_banks_20[209] = 32'h00000000;
assign filter_banks_20[210] = 32'h00000000;
assign filter_banks_20[211] = 32'h00000000;
assign filter_banks_20[212] = 32'h00000000;
assign filter_banks_20[213] = 32'h00000000;
assign filter_banks_20[214] = 32'h00000000;
assign filter_banks_20[215] = 32'h00000000;
assign filter_banks_20[216] = 32'h00000000;
assign filter_banks_20[217] = 32'h00000000;
assign filter_banks_20[218] = 32'h00000000;
assign filter_banks_20[219] = 32'h00000000;
assign filter_banks_20[220] = 32'h00000000;
assign filter_banks_20[221] = 32'h00000000;
assign filter_banks_20[222] = 32'h00000000;
assign filter_banks_20[223] = 32'h00000000;
assign filter_banks_20[224] = 32'h00000000;
assign filter_banks_20[225] = 32'h00000000;
assign filter_banks_20[226] = 32'h00000000;
assign filter_banks_20[227] = 32'h00000000;
assign filter_banks_20[228] = 32'h00000000;
assign filter_banks_20[229] = 32'h00000000;
assign filter_banks_20[230] = 32'h00000000;
assign filter_banks_20[231] = 32'h00000000;
assign filter_banks_20[232] = 32'h00000000;
assign filter_banks_20[233] = 32'h00000000;
assign filter_banks_20[234] = 32'h00000000;
assign filter_banks_20[235] = 32'h00000000;
assign filter_banks_20[236] = 32'h00000000;
assign filter_banks_20[237] = 32'h00000000;
assign filter_banks_20[238] = 32'h00000000;
assign filter_banks_20[239] = 32'h00000000;
assign filter_banks_20[240] = 32'h00000000;
assign filter_banks_20[241] = 32'h00000000;
assign filter_banks_20[242] = 32'h00000000;
assign filter_banks_20[243] = 32'h00000000;
assign filter_banks_20[244] = 32'h00000000;
assign filter_banks_20[245] = 32'h00000000;
assign filter_banks_20[246] = 32'h00000000;
assign filter_banks_20[247] = 32'h00000000;
assign filter_banks_20[248] = 32'h00000000;
assign filter_banks_20[249] = 32'h00000000;
assign filter_banks_20[250] = 32'h00000000;
assign filter_banks_20[251] = 32'h00000000;
assign filter_banks_20[252] = 32'h00000000;
assign filter_banks_20[253] = 32'h00000000;
assign filter_banks_20[254] = 32'h00000000;
assign filter_banks_20[255] = 32'h00000000;
assign filter_banks_20[256] = 32'h00000000;
assign filter_banks_21[0] = 32'h00000000;
assign filter_banks_21[1] = 32'h00000000;
assign filter_banks_21[2] = 32'h00000000;
assign filter_banks_21[3] = 32'h00000000;
assign filter_banks_21[4] = 32'h00000000;
assign filter_banks_21[5] = 32'h00000000;
assign filter_banks_21[6] = 32'h00000000;
assign filter_banks_21[7] = 32'h00000000;
assign filter_banks_21[8] = 32'h00000000;
assign filter_banks_21[9] = 32'h00000000;
assign filter_banks_21[10] = 32'h00000000;
assign filter_banks_21[11] = 32'h00000000;
assign filter_banks_21[12] = 32'h00000000;
assign filter_banks_21[13] = 32'h00000000;
assign filter_banks_21[14] = 32'h00000000;
assign filter_banks_21[15] = 32'h00000000;
assign filter_banks_21[16] = 32'h00000000;
assign filter_banks_21[17] = 32'h00000000;
assign filter_banks_21[18] = 32'h00000000;
assign filter_banks_21[19] = 32'h00000000;
assign filter_banks_21[20] = 32'h00000000;
assign filter_banks_21[21] = 32'h00000000;
assign filter_banks_21[22] = 32'h00000000;
assign filter_banks_21[23] = 32'h00000000;
assign filter_banks_21[24] = 32'h00000000;
assign filter_banks_21[25] = 32'h00000000;
assign filter_banks_21[26] = 32'h00000000;
assign filter_banks_21[27] = 32'h00000000;
assign filter_banks_21[28] = 32'h00000000;
assign filter_banks_21[29] = 32'h00000000;
assign filter_banks_21[30] = 32'h00000000;
assign filter_banks_21[31] = 32'h00000000;
assign filter_banks_21[32] = 32'h00000000;
assign filter_banks_21[33] = 32'h00000000;
assign filter_banks_21[34] = 32'h00000000;
assign filter_banks_21[35] = 32'h00000000;
assign filter_banks_21[36] = 32'h00000000;
assign filter_banks_21[37] = 32'h00000000;
assign filter_banks_21[38] = 32'h00000000;
assign filter_banks_21[39] = 32'h00000000;
assign filter_banks_21[40] = 32'h00000000;
assign filter_banks_21[41] = 32'h00000000;
assign filter_banks_21[42] = 32'h00000000;
assign filter_banks_21[43] = 32'h00000000;
assign filter_banks_21[44] = 32'h00000000;
assign filter_banks_21[45] = 32'h00000000;
assign filter_banks_21[46] = 32'h00000000;
assign filter_banks_21[47] = 32'h00000000;
assign filter_banks_21[48] = 32'h00000000;
assign filter_banks_21[49] = 32'h00000000;
assign filter_banks_21[50] = 32'h00000000;
assign filter_banks_21[51] = 32'h00000000;
assign filter_banks_21[52] = 32'h00000000;
assign filter_banks_21[53] = 32'h00000000;
assign filter_banks_21[54] = 32'h00000000;
assign filter_banks_21[55] = 32'h00000000;
assign filter_banks_21[56] = 32'h00000000;
assign filter_banks_21[57] = 32'h00000000;
assign filter_banks_21[58] = 32'h00000000;
assign filter_banks_21[59] = 32'h00000000;
assign filter_banks_21[60] = 32'h00000000;
assign filter_banks_21[61] = 32'h00000000;
assign filter_banks_21[62] = 32'h00000000;
assign filter_banks_21[63] = 32'h00000000;
assign filter_banks_21[64] = 32'h00000000;
assign filter_banks_21[65] = 32'h00000000;
assign filter_banks_21[66] = 32'h00000000;
assign filter_banks_21[67] = 32'h00000000;
assign filter_banks_21[68] = 32'h00000000;
assign filter_banks_21[69] = 32'h00000000;
assign filter_banks_21[70] = 32'h00000000;
assign filter_banks_21[71] = 32'h00000000;
assign filter_banks_21[72] = 32'h00000000;
assign filter_banks_21[73] = 32'h00000000;
assign filter_banks_21[74] = 32'h00000000;
assign filter_banks_21[75] = 32'h00000000;
assign filter_banks_21[76] = 32'h00000000;
assign filter_banks_21[77] = 32'h00000000;
assign filter_banks_21[78] = 32'h00000000;
assign filter_banks_21[79] = 32'h00000000;
assign filter_banks_21[80] = 32'h00000000;
assign filter_banks_21[81] = 32'h00000000;
assign filter_banks_21[82] = 32'h00000000;
assign filter_banks_21[83] = 32'h00000000;
assign filter_banks_21[84] = 32'h00000000;
assign filter_banks_21[85] = 32'h00000000;
assign filter_banks_21[86] = 32'h00000000;
assign filter_banks_21[87] = 32'h00000000;
assign filter_banks_21[88] = 32'h00000000;
assign filter_banks_21[89] = 32'h00000000;
assign filter_banks_21[90] = 32'h00000000;
assign filter_banks_21[91] = 32'h00000000;
assign filter_banks_21[92] = 32'h00000000;
assign filter_banks_21[93] = 32'h00000000;
assign filter_banks_21[94] = 32'h00000000;
assign filter_banks_21[95] = 32'h00000000;
assign filter_banks_21[96] = 32'h00000000;
assign filter_banks_21[97] = 32'h00000000;
assign filter_banks_21[98] = 32'h00000000;
assign filter_banks_21[99] = 32'h00000000;
assign filter_banks_21[100] = 32'h00000000;
assign filter_banks_21[101] = 32'h00000000;
assign filter_banks_21[102] = 32'h00000000;
assign filter_banks_21[103] = 32'h00000000;
assign filter_banks_21[104] = 32'h00000000;
assign filter_banks_21[105] = 32'h00000000;
assign filter_banks_21[106] = 32'h00000000;
assign filter_banks_21[107] = 32'h00000000;
assign filter_banks_21[108] = 32'h00000000;
assign filter_banks_21[109] = 32'h00000000;
assign filter_banks_21[110] = 32'h00000000;
assign filter_banks_21[111] = 32'h00000000;
assign filter_banks_21[112] = 32'h00000000;
assign filter_banks_21[113] = 32'h00000000;
assign filter_banks_21[114] = 32'h00000000;
assign filter_banks_21[115] = 32'h00000000;
assign filter_banks_21[116] = 32'h00000000;
assign filter_banks_21[117] = 32'h00000000;
assign filter_banks_21[118] = 32'h00000000;
assign filter_banks_21[119] = 32'h00000000;
assign filter_banks_21[120] = 32'h00000000;
assign filter_banks_21[121] = 32'h00000000;
assign filter_banks_21[122] = 32'h00000000;
assign filter_banks_21[123] = 32'h3d924925;
assign filter_banks_21[124] = 32'h3e124925;
assign filter_banks_21[125] = 32'h3e5b6db7;
assign filter_banks_21[126] = 32'h3e924925;
assign filter_banks_21[127] = 32'h3eb6db6e;
assign filter_banks_21[128] = 32'h3edb6db7;
assign filter_banks_21[129] = 32'h3f000000;
assign filter_banks_21[130] = 32'h3f124925;
assign filter_banks_21[131] = 32'h3f249249;
assign filter_banks_21[132] = 32'h3f36db6e;
assign filter_banks_21[133] = 32'h3f492492;
assign filter_banks_21[134] = 32'h3f5b6db7;
assign filter_banks_21[135] = 32'h3f6db6db;
assign filter_banks_21[136] = 32'h3f800000;
assign filter_banks_21[137] = 32'h3f700000;
assign filter_banks_21[138] = 32'h3f600000;
assign filter_banks_21[139] = 32'h3f500000;
assign filter_banks_21[140] = 32'h3f400000;
assign filter_banks_21[141] = 32'h3f300000;
assign filter_banks_21[142] = 32'h3f200000;
assign filter_banks_21[143] = 32'h3f100000;
assign filter_banks_21[144] = 32'h3f000000;
assign filter_banks_21[145] = 32'h3ee00000;
assign filter_banks_21[146] = 32'h3ec00000;
assign filter_banks_21[147] = 32'h3ea00000;
assign filter_banks_21[148] = 32'h3e800000;
assign filter_banks_21[149] = 32'h3e400000;
assign filter_banks_21[150] = 32'h3e000000;
assign filter_banks_21[151] = 32'h3d800000;
assign filter_banks_21[152] = 32'h00000000;
assign filter_banks_21[153] = 32'h00000000;
assign filter_banks_21[154] = 32'h00000000;
assign filter_banks_21[155] = 32'h00000000;
assign filter_banks_21[156] = 32'h00000000;
assign filter_banks_21[157] = 32'h00000000;
assign filter_banks_21[158] = 32'h00000000;
assign filter_banks_21[159] = 32'h00000000;
assign filter_banks_21[160] = 32'h00000000;
assign filter_banks_21[161] = 32'h00000000;
assign filter_banks_21[162] = 32'h00000000;
assign filter_banks_21[163] = 32'h00000000;
assign filter_banks_21[164] = 32'h00000000;
assign filter_banks_21[165] = 32'h00000000;
assign filter_banks_21[166] = 32'h00000000;
assign filter_banks_21[167] = 32'h00000000;
assign filter_banks_21[168] = 32'h00000000;
assign filter_banks_21[169] = 32'h00000000;
assign filter_banks_21[170] = 32'h00000000;
assign filter_banks_21[171] = 32'h00000000;
assign filter_banks_21[172] = 32'h00000000;
assign filter_banks_21[173] = 32'h00000000;
assign filter_banks_21[174] = 32'h00000000;
assign filter_banks_21[175] = 32'h00000000;
assign filter_banks_21[176] = 32'h00000000;
assign filter_banks_21[177] = 32'h00000000;
assign filter_banks_21[178] = 32'h00000000;
assign filter_banks_21[179] = 32'h00000000;
assign filter_banks_21[180] = 32'h00000000;
assign filter_banks_21[181] = 32'h00000000;
assign filter_banks_21[182] = 32'h00000000;
assign filter_banks_21[183] = 32'h00000000;
assign filter_banks_21[184] = 32'h00000000;
assign filter_banks_21[185] = 32'h00000000;
assign filter_banks_21[186] = 32'h00000000;
assign filter_banks_21[187] = 32'h00000000;
assign filter_banks_21[188] = 32'h00000000;
assign filter_banks_21[189] = 32'h00000000;
assign filter_banks_21[190] = 32'h00000000;
assign filter_banks_21[191] = 32'h00000000;
assign filter_banks_21[192] = 32'h00000000;
assign filter_banks_21[193] = 32'h00000000;
assign filter_banks_21[194] = 32'h00000000;
assign filter_banks_21[195] = 32'h00000000;
assign filter_banks_21[196] = 32'h00000000;
assign filter_banks_21[197] = 32'h00000000;
assign filter_banks_21[198] = 32'h00000000;
assign filter_banks_21[199] = 32'h00000000;
assign filter_banks_21[200] = 32'h00000000;
assign filter_banks_21[201] = 32'h00000000;
assign filter_banks_21[202] = 32'h00000000;
assign filter_banks_21[203] = 32'h00000000;
assign filter_banks_21[204] = 32'h00000000;
assign filter_banks_21[205] = 32'h00000000;
assign filter_banks_21[206] = 32'h00000000;
assign filter_banks_21[207] = 32'h00000000;
assign filter_banks_21[208] = 32'h00000000;
assign filter_banks_21[209] = 32'h00000000;
assign filter_banks_21[210] = 32'h00000000;
assign filter_banks_21[211] = 32'h00000000;
assign filter_banks_21[212] = 32'h00000000;
assign filter_banks_21[213] = 32'h00000000;
assign filter_banks_21[214] = 32'h00000000;
assign filter_banks_21[215] = 32'h00000000;
assign filter_banks_21[216] = 32'h00000000;
assign filter_banks_21[217] = 32'h00000000;
assign filter_banks_21[218] = 32'h00000000;
assign filter_banks_21[219] = 32'h00000000;
assign filter_banks_21[220] = 32'h00000000;
assign filter_banks_21[221] = 32'h00000000;
assign filter_banks_21[222] = 32'h00000000;
assign filter_banks_21[223] = 32'h00000000;
assign filter_banks_21[224] = 32'h00000000;
assign filter_banks_21[225] = 32'h00000000;
assign filter_banks_21[226] = 32'h00000000;
assign filter_banks_21[227] = 32'h00000000;
assign filter_banks_21[228] = 32'h00000000;
assign filter_banks_21[229] = 32'h00000000;
assign filter_banks_21[230] = 32'h00000000;
assign filter_banks_21[231] = 32'h00000000;
assign filter_banks_21[232] = 32'h00000000;
assign filter_banks_21[233] = 32'h00000000;
assign filter_banks_21[234] = 32'h00000000;
assign filter_banks_21[235] = 32'h00000000;
assign filter_banks_21[236] = 32'h00000000;
assign filter_banks_21[237] = 32'h00000000;
assign filter_banks_21[238] = 32'h00000000;
assign filter_banks_21[239] = 32'h00000000;
assign filter_banks_21[240] = 32'h00000000;
assign filter_banks_21[241] = 32'h00000000;
assign filter_banks_21[242] = 32'h00000000;
assign filter_banks_21[243] = 32'h00000000;
assign filter_banks_21[244] = 32'h00000000;
assign filter_banks_21[245] = 32'h00000000;
assign filter_banks_21[246] = 32'h00000000;
assign filter_banks_21[247] = 32'h00000000;
assign filter_banks_21[248] = 32'h00000000;
assign filter_banks_21[249] = 32'h00000000;
assign filter_banks_21[250] = 32'h00000000;
assign filter_banks_21[251] = 32'h00000000;
assign filter_banks_21[252] = 32'h00000000;
assign filter_banks_21[253] = 32'h00000000;
assign filter_banks_21[254] = 32'h00000000;
assign filter_banks_21[255] = 32'h00000000;
assign filter_banks_21[256] = 32'h00000000;
assign filter_banks_22[0] = 32'h00000000;
assign filter_banks_22[1] = 32'h00000000;
assign filter_banks_22[2] = 32'h00000000;
assign filter_banks_22[3] = 32'h00000000;
assign filter_banks_22[4] = 32'h00000000;
assign filter_banks_22[5] = 32'h00000000;
assign filter_banks_22[6] = 32'h00000000;
assign filter_banks_22[7] = 32'h00000000;
assign filter_banks_22[8] = 32'h00000000;
assign filter_banks_22[9] = 32'h00000000;
assign filter_banks_22[10] = 32'h00000000;
assign filter_banks_22[11] = 32'h00000000;
assign filter_banks_22[12] = 32'h00000000;
assign filter_banks_22[13] = 32'h00000000;
assign filter_banks_22[14] = 32'h00000000;
assign filter_banks_22[15] = 32'h00000000;
assign filter_banks_22[16] = 32'h00000000;
assign filter_banks_22[17] = 32'h00000000;
assign filter_banks_22[18] = 32'h00000000;
assign filter_banks_22[19] = 32'h00000000;
assign filter_banks_22[20] = 32'h00000000;
assign filter_banks_22[21] = 32'h00000000;
assign filter_banks_22[22] = 32'h00000000;
assign filter_banks_22[23] = 32'h00000000;
assign filter_banks_22[24] = 32'h00000000;
assign filter_banks_22[25] = 32'h00000000;
assign filter_banks_22[26] = 32'h00000000;
assign filter_banks_22[27] = 32'h00000000;
assign filter_banks_22[28] = 32'h00000000;
assign filter_banks_22[29] = 32'h00000000;
assign filter_banks_22[30] = 32'h00000000;
assign filter_banks_22[31] = 32'h00000000;
assign filter_banks_22[32] = 32'h00000000;
assign filter_banks_22[33] = 32'h00000000;
assign filter_banks_22[34] = 32'h00000000;
assign filter_banks_22[35] = 32'h00000000;
assign filter_banks_22[36] = 32'h00000000;
assign filter_banks_22[37] = 32'h00000000;
assign filter_banks_22[38] = 32'h00000000;
assign filter_banks_22[39] = 32'h00000000;
assign filter_banks_22[40] = 32'h00000000;
assign filter_banks_22[41] = 32'h00000000;
assign filter_banks_22[42] = 32'h00000000;
assign filter_banks_22[43] = 32'h00000000;
assign filter_banks_22[44] = 32'h00000000;
assign filter_banks_22[45] = 32'h00000000;
assign filter_banks_22[46] = 32'h00000000;
assign filter_banks_22[47] = 32'h00000000;
assign filter_banks_22[48] = 32'h00000000;
assign filter_banks_22[49] = 32'h00000000;
assign filter_banks_22[50] = 32'h00000000;
assign filter_banks_22[51] = 32'h00000000;
assign filter_banks_22[52] = 32'h00000000;
assign filter_banks_22[53] = 32'h00000000;
assign filter_banks_22[54] = 32'h00000000;
assign filter_banks_22[55] = 32'h00000000;
assign filter_banks_22[56] = 32'h00000000;
assign filter_banks_22[57] = 32'h00000000;
assign filter_banks_22[58] = 32'h00000000;
assign filter_banks_22[59] = 32'h00000000;
assign filter_banks_22[60] = 32'h00000000;
assign filter_banks_22[61] = 32'h00000000;
assign filter_banks_22[62] = 32'h00000000;
assign filter_banks_22[63] = 32'h00000000;
assign filter_banks_22[64] = 32'h00000000;
assign filter_banks_22[65] = 32'h00000000;
assign filter_banks_22[66] = 32'h00000000;
assign filter_banks_22[67] = 32'h00000000;
assign filter_banks_22[68] = 32'h00000000;
assign filter_banks_22[69] = 32'h00000000;
assign filter_banks_22[70] = 32'h00000000;
assign filter_banks_22[71] = 32'h00000000;
assign filter_banks_22[72] = 32'h00000000;
assign filter_banks_22[73] = 32'h00000000;
assign filter_banks_22[74] = 32'h00000000;
assign filter_banks_22[75] = 32'h00000000;
assign filter_banks_22[76] = 32'h00000000;
assign filter_banks_22[77] = 32'h00000000;
assign filter_banks_22[78] = 32'h00000000;
assign filter_banks_22[79] = 32'h00000000;
assign filter_banks_22[80] = 32'h00000000;
assign filter_banks_22[81] = 32'h00000000;
assign filter_banks_22[82] = 32'h00000000;
assign filter_banks_22[83] = 32'h00000000;
assign filter_banks_22[84] = 32'h00000000;
assign filter_banks_22[85] = 32'h00000000;
assign filter_banks_22[86] = 32'h00000000;
assign filter_banks_22[87] = 32'h00000000;
assign filter_banks_22[88] = 32'h00000000;
assign filter_banks_22[89] = 32'h00000000;
assign filter_banks_22[90] = 32'h00000000;
assign filter_banks_22[91] = 32'h00000000;
assign filter_banks_22[92] = 32'h00000000;
assign filter_banks_22[93] = 32'h00000000;
assign filter_banks_22[94] = 32'h00000000;
assign filter_banks_22[95] = 32'h00000000;
assign filter_banks_22[96] = 32'h00000000;
assign filter_banks_22[97] = 32'h00000000;
assign filter_banks_22[98] = 32'h00000000;
assign filter_banks_22[99] = 32'h00000000;
assign filter_banks_22[100] = 32'h00000000;
assign filter_banks_22[101] = 32'h00000000;
assign filter_banks_22[102] = 32'h00000000;
assign filter_banks_22[103] = 32'h00000000;
assign filter_banks_22[104] = 32'h00000000;
assign filter_banks_22[105] = 32'h00000000;
assign filter_banks_22[106] = 32'h00000000;
assign filter_banks_22[107] = 32'h00000000;
assign filter_banks_22[108] = 32'h00000000;
assign filter_banks_22[109] = 32'h00000000;
assign filter_banks_22[110] = 32'h00000000;
assign filter_banks_22[111] = 32'h00000000;
assign filter_banks_22[112] = 32'h00000000;
assign filter_banks_22[113] = 32'h00000000;
assign filter_banks_22[114] = 32'h00000000;
assign filter_banks_22[115] = 32'h00000000;
assign filter_banks_22[116] = 32'h00000000;
assign filter_banks_22[117] = 32'h00000000;
assign filter_banks_22[118] = 32'h00000000;
assign filter_banks_22[119] = 32'h00000000;
assign filter_banks_22[120] = 32'h00000000;
assign filter_banks_22[121] = 32'h00000000;
assign filter_banks_22[122] = 32'h00000000;
assign filter_banks_22[123] = 32'h00000000;
assign filter_banks_22[124] = 32'h00000000;
assign filter_banks_22[125] = 32'h00000000;
assign filter_banks_22[126] = 32'h00000000;
assign filter_banks_22[127] = 32'h00000000;
assign filter_banks_22[128] = 32'h00000000;
assign filter_banks_22[129] = 32'h00000000;
assign filter_banks_22[130] = 32'h00000000;
assign filter_banks_22[131] = 32'h00000000;
assign filter_banks_22[132] = 32'h00000000;
assign filter_banks_22[133] = 32'h00000000;
assign filter_banks_22[134] = 32'h00000000;
assign filter_banks_22[135] = 32'h00000000;
assign filter_banks_22[136] = 32'h00000000;
assign filter_banks_22[137] = 32'h3d800000;
assign filter_banks_22[138] = 32'h3e000000;
assign filter_banks_22[139] = 32'h3e400000;
assign filter_banks_22[140] = 32'h3e800000;
assign filter_banks_22[141] = 32'h3ea00000;
assign filter_banks_22[142] = 32'h3ec00000;
assign filter_banks_22[143] = 32'h3ee00000;
assign filter_banks_22[144] = 32'h3f000000;
assign filter_banks_22[145] = 32'h3f100000;
assign filter_banks_22[146] = 32'h3f200000;
assign filter_banks_22[147] = 32'h3f300000;
assign filter_banks_22[148] = 32'h3f400000;
assign filter_banks_22[149] = 32'h3f500000;
assign filter_banks_22[150] = 32'h3f600000;
assign filter_banks_22[151] = 32'h3f700000;
assign filter_banks_22[152] = 32'h3f800000;
assign filter_banks_22[153] = 32'h3f70f0f1;
assign filter_banks_22[154] = 32'h3f61e1e2;
assign filter_banks_22[155] = 32'h3f52d2d3;
assign filter_banks_22[156] = 32'h3f43c3c4;
assign filter_banks_22[157] = 32'h3f34b4b5;
assign filter_banks_22[158] = 32'h3f25a5a6;
assign filter_banks_22[159] = 32'h3f169697;
assign filter_banks_22[160] = 32'h3f078788;
assign filter_banks_22[161] = 32'h3ef0f0f1;
assign filter_banks_22[162] = 32'h3ed2d2d3;
assign filter_banks_22[163] = 32'h3eb4b4b5;
assign filter_banks_22[164] = 32'h3e969697;
assign filter_banks_22[165] = 32'h3e70f0f1;
assign filter_banks_22[166] = 32'h3e34b4b5;
assign filter_banks_22[167] = 32'h3df0f0f1;
assign filter_banks_22[168] = 32'h3d70f0f1;
assign filter_banks_22[169] = 32'h00000000;
assign filter_banks_22[170] = 32'h00000000;
assign filter_banks_22[171] = 32'h00000000;
assign filter_banks_22[172] = 32'h00000000;
assign filter_banks_22[173] = 32'h00000000;
assign filter_banks_22[174] = 32'h00000000;
assign filter_banks_22[175] = 32'h00000000;
assign filter_banks_22[176] = 32'h00000000;
assign filter_banks_22[177] = 32'h00000000;
assign filter_banks_22[178] = 32'h00000000;
assign filter_banks_22[179] = 32'h00000000;
assign filter_banks_22[180] = 32'h00000000;
assign filter_banks_22[181] = 32'h00000000;
assign filter_banks_22[182] = 32'h00000000;
assign filter_banks_22[183] = 32'h00000000;
assign filter_banks_22[184] = 32'h00000000;
assign filter_banks_22[185] = 32'h00000000;
assign filter_banks_22[186] = 32'h00000000;
assign filter_banks_22[187] = 32'h00000000;
assign filter_banks_22[188] = 32'h00000000;
assign filter_banks_22[189] = 32'h00000000;
assign filter_banks_22[190] = 32'h00000000;
assign filter_banks_22[191] = 32'h00000000;
assign filter_banks_22[192] = 32'h00000000;
assign filter_banks_22[193] = 32'h00000000;
assign filter_banks_22[194] = 32'h00000000;
assign filter_banks_22[195] = 32'h00000000;
assign filter_banks_22[196] = 32'h00000000;
assign filter_banks_22[197] = 32'h00000000;
assign filter_banks_22[198] = 32'h00000000;
assign filter_banks_22[199] = 32'h00000000;
assign filter_banks_22[200] = 32'h00000000;
assign filter_banks_22[201] = 32'h00000000;
assign filter_banks_22[202] = 32'h00000000;
assign filter_banks_22[203] = 32'h00000000;
assign filter_banks_22[204] = 32'h00000000;
assign filter_banks_22[205] = 32'h00000000;
assign filter_banks_22[206] = 32'h00000000;
assign filter_banks_22[207] = 32'h00000000;
assign filter_banks_22[208] = 32'h00000000;
assign filter_banks_22[209] = 32'h00000000;
assign filter_banks_22[210] = 32'h00000000;
assign filter_banks_22[211] = 32'h00000000;
assign filter_banks_22[212] = 32'h00000000;
assign filter_banks_22[213] = 32'h00000000;
assign filter_banks_22[214] = 32'h00000000;
assign filter_banks_22[215] = 32'h00000000;
assign filter_banks_22[216] = 32'h00000000;
assign filter_banks_22[217] = 32'h00000000;
assign filter_banks_22[218] = 32'h00000000;
assign filter_banks_22[219] = 32'h00000000;
assign filter_banks_22[220] = 32'h00000000;
assign filter_banks_22[221] = 32'h00000000;
assign filter_banks_22[222] = 32'h00000000;
assign filter_banks_22[223] = 32'h00000000;
assign filter_banks_22[224] = 32'h00000000;
assign filter_banks_22[225] = 32'h00000000;
assign filter_banks_22[226] = 32'h00000000;
assign filter_banks_22[227] = 32'h00000000;
assign filter_banks_22[228] = 32'h00000000;
assign filter_banks_22[229] = 32'h00000000;
assign filter_banks_22[230] = 32'h00000000;
assign filter_banks_22[231] = 32'h00000000;
assign filter_banks_22[232] = 32'h00000000;
assign filter_banks_22[233] = 32'h00000000;
assign filter_banks_22[234] = 32'h00000000;
assign filter_banks_22[235] = 32'h00000000;
assign filter_banks_22[236] = 32'h00000000;
assign filter_banks_22[237] = 32'h00000000;
assign filter_banks_22[238] = 32'h00000000;
assign filter_banks_22[239] = 32'h00000000;
assign filter_banks_22[240] = 32'h00000000;
assign filter_banks_22[241] = 32'h00000000;
assign filter_banks_22[242] = 32'h00000000;
assign filter_banks_22[243] = 32'h00000000;
assign filter_banks_22[244] = 32'h00000000;
assign filter_banks_22[245] = 32'h00000000;
assign filter_banks_22[246] = 32'h00000000;
assign filter_banks_22[247] = 32'h00000000;
assign filter_banks_22[248] = 32'h00000000;
assign filter_banks_22[249] = 32'h00000000;
assign filter_banks_22[250] = 32'h00000000;
assign filter_banks_22[251] = 32'h00000000;
assign filter_banks_22[252] = 32'h00000000;
assign filter_banks_22[253] = 32'h00000000;
assign filter_banks_22[254] = 32'h00000000;
assign filter_banks_22[255] = 32'h00000000;
assign filter_banks_22[256] = 32'h00000000;
assign filter_banks_23[0] = 32'h00000000;
assign filter_banks_23[1] = 32'h00000000;
assign filter_banks_23[2] = 32'h00000000;
assign filter_banks_23[3] = 32'h00000000;
assign filter_banks_23[4] = 32'h00000000;
assign filter_banks_23[5] = 32'h00000000;
assign filter_banks_23[6] = 32'h00000000;
assign filter_banks_23[7] = 32'h00000000;
assign filter_banks_23[8] = 32'h00000000;
assign filter_banks_23[9] = 32'h00000000;
assign filter_banks_23[10] = 32'h00000000;
assign filter_banks_23[11] = 32'h00000000;
assign filter_banks_23[12] = 32'h00000000;
assign filter_banks_23[13] = 32'h00000000;
assign filter_banks_23[14] = 32'h00000000;
assign filter_banks_23[15] = 32'h00000000;
assign filter_banks_23[16] = 32'h00000000;
assign filter_banks_23[17] = 32'h00000000;
assign filter_banks_23[18] = 32'h00000000;
assign filter_banks_23[19] = 32'h00000000;
assign filter_banks_23[20] = 32'h00000000;
assign filter_banks_23[21] = 32'h00000000;
assign filter_banks_23[22] = 32'h00000000;
assign filter_banks_23[23] = 32'h00000000;
assign filter_banks_23[24] = 32'h00000000;
assign filter_banks_23[25] = 32'h00000000;
assign filter_banks_23[26] = 32'h00000000;
assign filter_banks_23[27] = 32'h00000000;
assign filter_banks_23[28] = 32'h00000000;
assign filter_banks_23[29] = 32'h00000000;
assign filter_banks_23[30] = 32'h00000000;
assign filter_banks_23[31] = 32'h00000000;
assign filter_banks_23[32] = 32'h00000000;
assign filter_banks_23[33] = 32'h00000000;
assign filter_banks_23[34] = 32'h00000000;
assign filter_banks_23[35] = 32'h00000000;
assign filter_banks_23[36] = 32'h00000000;
assign filter_banks_23[37] = 32'h00000000;
assign filter_banks_23[38] = 32'h00000000;
assign filter_banks_23[39] = 32'h00000000;
assign filter_banks_23[40] = 32'h00000000;
assign filter_banks_23[41] = 32'h00000000;
assign filter_banks_23[42] = 32'h00000000;
assign filter_banks_23[43] = 32'h00000000;
assign filter_banks_23[44] = 32'h00000000;
assign filter_banks_23[45] = 32'h00000000;
assign filter_banks_23[46] = 32'h00000000;
assign filter_banks_23[47] = 32'h00000000;
assign filter_banks_23[48] = 32'h00000000;
assign filter_banks_23[49] = 32'h00000000;
assign filter_banks_23[50] = 32'h00000000;
assign filter_banks_23[51] = 32'h00000000;
assign filter_banks_23[52] = 32'h00000000;
assign filter_banks_23[53] = 32'h00000000;
assign filter_banks_23[54] = 32'h00000000;
assign filter_banks_23[55] = 32'h00000000;
assign filter_banks_23[56] = 32'h00000000;
assign filter_banks_23[57] = 32'h00000000;
assign filter_banks_23[58] = 32'h00000000;
assign filter_banks_23[59] = 32'h00000000;
assign filter_banks_23[60] = 32'h00000000;
assign filter_banks_23[61] = 32'h00000000;
assign filter_banks_23[62] = 32'h00000000;
assign filter_banks_23[63] = 32'h00000000;
assign filter_banks_23[64] = 32'h00000000;
assign filter_banks_23[65] = 32'h00000000;
assign filter_banks_23[66] = 32'h00000000;
assign filter_banks_23[67] = 32'h00000000;
assign filter_banks_23[68] = 32'h00000000;
assign filter_banks_23[69] = 32'h00000000;
assign filter_banks_23[70] = 32'h00000000;
assign filter_banks_23[71] = 32'h00000000;
assign filter_banks_23[72] = 32'h00000000;
assign filter_banks_23[73] = 32'h00000000;
assign filter_banks_23[74] = 32'h00000000;
assign filter_banks_23[75] = 32'h00000000;
assign filter_banks_23[76] = 32'h00000000;
assign filter_banks_23[77] = 32'h00000000;
assign filter_banks_23[78] = 32'h00000000;
assign filter_banks_23[79] = 32'h00000000;
assign filter_banks_23[80] = 32'h00000000;
assign filter_banks_23[81] = 32'h00000000;
assign filter_banks_23[82] = 32'h00000000;
assign filter_banks_23[83] = 32'h00000000;
assign filter_banks_23[84] = 32'h00000000;
assign filter_banks_23[85] = 32'h00000000;
assign filter_banks_23[86] = 32'h00000000;
assign filter_banks_23[87] = 32'h00000000;
assign filter_banks_23[88] = 32'h00000000;
assign filter_banks_23[89] = 32'h00000000;
assign filter_banks_23[90] = 32'h00000000;
assign filter_banks_23[91] = 32'h00000000;
assign filter_banks_23[92] = 32'h00000000;
assign filter_banks_23[93] = 32'h00000000;
assign filter_banks_23[94] = 32'h00000000;
assign filter_banks_23[95] = 32'h00000000;
assign filter_banks_23[96] = 32'h00000000;
assign filter_banks_23[97] = 32'h00000000;
assign filter_banks_23[98] = 32'h00000000;
assign filter_banks_23[99] = 32'h00000000;
assign filter_banks_23[100] = 32'h00000000;
assign filter_banks_23[101] = 32'h00000000;
assign filter_banks_23[102] = 32'h00000000;
assign filter_banks_23[103] = 32'h00000000;
assign filter_banks_23[104] = 32'h00000000;
assign filter_banks_23[105] = 32'h00000000;
assign filter_banks_23[106] = 32'h00000000;
assign filter_banks_23[107] = 32'h00000000;
assign filter_banks_23[108] = 32'h00000000;
assign filter_banks_23[109] = 32'h00000000;
assign filter_banks_23[110] = 32'h00000000;
assign filter_banks_23[111] = 32'h00000000;
assign filter_banks_23[112] = 32'h00000000;
assign filter_banks_23[113] = 32'h00000000;
assign filter_banks_23[114] = 32'h00000000;
assign filter_banks_23[115] = 32'h00000000;
assign filter_banks_23[116] = 32'h00000000;
assign filter_banks_23[117] = 32'h00000000;
assign filter_banks_23[118] = 32'h00000000;
assign filter_banks_23[119] = 32'h00000000;
assign filter_banks_23[120] = 32'h00000000;
assign filter_banks_23[121] = 32'h00000000;
assign filter_banks_23[122] = 32'h00000000;
assign filter_banks_23[123] = 32'h00000000;
assign filter_banks_23[124] = 32'h00000000;
assign filter_banks_23[125] = 32'h00000000;
assign filter_banks_23[126] = 32'h00000000;
assign filter_banks_23[127] = 32'h00000000;
assign filter_banks_23[128] = 32'h00000000;
assign filter_banks_23[129] = 32'h00000000;
assign filter_banks_23[130] = 32'h00000000;
assign filter_banks_23[131] = 32'h00000000;
assign filter_banks_23[132] = 32'h00000000;
assign filter_banks_23[133] = 32'h00000000;
assign filter_banks_23[134] = 32'h00000000;
assign filter_banks_23[135] = 32'h00000000;
assign filter_banks_23[136] = 32'h00000000;
assign filter_banks_23[137] = 32'h00000000;
assign filter_banks_23[138] = 32'h00000000;
assign filter_banks_23[139] = 32'h00000000;
assign filter_banks_23[140] = 32'h00000000;
assign filter_banks_23[141] = 32'h00000000;
assign filter_banks_23[142] = 32'h00000000;
assign filter_banks_23[143] = 32'h00000000;
assign filter_banks_23[144] = 32'h00000000;
assign filter_banks_23[145] = 32'h00000000;
assign filter_banks_23[146] = 32'h00000000;
assign filter_banks_23[147] = 32'h00000000;
assign filter_banks_23[148] = 32'h00000000;
assign filter_banks_23[149] = 32'h00000000;
assign filter_banks_23[150] = 32'h00000000;
assign filter_banks_23[151] = 32'h00000000;
assign filter_banks_23[152] = 32'h00000000;
assign filter_banks_23[153] = 32'h3d70f0f1;
assign filter_banks_23[154] = 32'h3df0f0f1;
assign filter_banks_23[155] = 32'h3e34b4b5;
assign filter_banks_23[156] = 32'h3e70f0f1;
assign filter_banks_23[157] = 32'h3e969697;
assign filter_banks_23[158] = 32'h3eb4b4b5;
assign filter_banks_23[159] = 32'h3ed2d2d3;
assign filter_banks_23[160] = 32'h3ef0f0f1;
assign filter_banks_23[161] = 32'h3f078788;
assign filter_banks_23[162] = 32'h3f169697;
assign filter_banks_23[163] = 32'h3f25a5a6;
assign filter_banks_23[164] = 32'h3f34b4b5;
assign filter_banks_23[165] = 32'h3f43c3c4;
assign filter_banks_23[166] = 32'h3f52d2d3;
assign filter_banks_23[167] = 32'h3f61e1e2;
assign filter_banks_23[168] = 32'h3f70f0f1;
assign filter_banks_23[169] = 32'h3f800000;
assign filter_banks_23[170] = 32'h3f7286bd;
assign filter_banks_23[171] = 32'h3f650d79;
assign filter_banks_23[172] = 32'h3f579436;
assign filter_banks_23[173] = 32'h3f4a1af3;
assign filter_banks_23[174] = 32'h3f3ca1af;
assign filter_banks_23[175] = 32'h3f2f286c;
assign filter_banks_23[176] = 32'h3f21af28;
assign filter_banks_23[177] = 32'h3f1435e5;
assign filter_banks_23[178] = 32'h3f06bca2;
assign filter_banks_23[179] = 32'h3ef286bd;
assign filter_banks_23[180] = 32'h3ed79436;
assign filter_banks_23[181] = 32'h3ebca1af;
assign filter_banks_23[182] = 32'h3ea1af28;
assign filter_banks_23[183] = 32'h3e86bca2;
assign filter_banks_23[184] = 32'h3e579436;
assign filter_banks_23[185] = 32'h3e21af28;
assign filter_banks_23[186] = 32'h3dd79436;
assign filter_banks_23[187] = 32'h3d579436;
assign filter_banks_23[188] = 32'h00000000;
assign filter_banks_23[189] = 32'h00000000;
assign filter_banks_23[190] = 32'h00000000;
assign filter_banks_23[191] = 32'h00000000;
assign filter_banks_23[192] = 32'h00000000;
assign filter_banks_23[193] = 32'h00000000;
assign filter_banks_23[194] = 32'h00000000;
assign filter_banks_23[195] = 32'h00000000;
assign filter_banks_23[196] = 32'h00000000;
assign filter_banks_23[197] = 32'h00000000;
assign filter_banks_23[198] = 32'h00000000;
assign filter_banks_23[199] = 32'h00000000;
assign filter_banks_23[200] = 32'h00000000;
assign filter_banks_23[201] = 32'h00000000;
assign filter_banks_23[202] = 32'h00000000;
assign filter_banks_23[203] = 32'h00000000;
assign filter_banks_23[204] = 32'h00000000;
assign filter_banks_23[205] = 32'h00000000;
assign filter_banks_23[206] = 32'h00000000;
assign filter_banks_23[207] = 32'h00000000;
assign filter_banks_23[208] = 32'h00000000;
assign filter_banks_23[209] = 32'h00000000;
assign filter_banks_23[210] = 32'h00000000;
assign filter_banks_23[211] = 32'h00000000;
assign filter_banks_23[212] = 32'h00000000;
assign filter_banks_23[213] = 32'h00000000;
assign filter_banks_23[214] = 32'h00000000;
assign filter_banks_23[215] = 32'h00000000;
assign filter_banks_23[216] = 32'h00000000;
assign filter_banks_23[217] = 32'h00000000;
assign filter_banks_23[218] = 32'h00000000;
assign filter_banks_23[219] = 32'h00000000;
assign filter_banks_23[220] = 32'h00000000;
assign filter_banks_23[221] = 32'h00000000;
assign filter_banks_23[222] = 32'h00000000;
assign filter_banks_23[223] = 32'h00000000;
assign filter_banks_23[224] = 32'h00000000;
assign filter_banks_23[225] = 32'h00000000;
assign filter_banks_23[226] = 32'h00000000;
assign filter_banks_23[227] = 32'h00000000;
assign filter_banks_23[228] = 32'h00000000;
assign filter_banks_23[229] = 32'h00000000;
assign filter_banks_23[230] = 32'h00000000;
assign filter_banks_23[231] = 32'h00000000;
assign filter_banks_23[232] = 32'h00000000;
assign filter_banks_23[233] = 32'h00000000;
assign filter_banks_23[234] = 32'h00000000;
assign filter_banks_23[235] = 32'h00000000;
assign filter_banks_23[236] = 32'h00000000;
assign filter_banks_23[237] = 32'h00000000;
assign filter_banks_23[238] = 32'h00000000;
assign filter_banks_23[239] = 32'h00000000;
assign filter_banks_23[240] = 32'h00000000;
assign filter_banks_23[241] = 32'h00000000;
assign filter_banks_23[242] = 32'h00000000;
assign filter_banks_23[243] = 32'h00000000;
assign filter_banks_23[244] = 32'h00000000;
assign filter_banks_23[245] = 32'h00000000;
assign filter_banks_23[246] = 32'h00000000;
assign filter_banks_23[247] = 32'h00000000;
assign filter_banks_23[248] = 32'h00000000;
assign filter_banks_23[249] = 32'h00000000;
assign filter_banks_23[250] = 32'h00000000;
assign filter_banks_23[251] = 32'h00000000;
assign filter_banks_23[252] = 32'h00000000;
assign filter_banks_23[253] = 32'h00000000;
assign filter_banks_23[254] = 32'h00000000;
assign filter_banks_23[255] = 32'h00000000;
assign filter_banks_23[256] = 32'h00000000;
assign filter_banks_24[0] = 32'h00000000;
assign filter_banks_24[1] = 32'h00000000;
assign filter_banks_24[2] = 32'h00000000;
assign filter_banks_24[3] = 32'h00000000;
assign filter_banks_24[4] = 32'h00000000;
assign filter_banks_24[5] = 32'h00000000;
assign filter_banks_24[6] = 32'h00000000;
assign filter_banks_24[7] = 32'h00000000;
assign filter_banks_24[8] = 32'h00000000;
assign filter_banks_24[9] = 32'h00000000;
assign filter_banks_24[10] = 32'h00000000;
assign filter_banks_24[11] = 32'h00000000;
assign filter_banks_24[12] = 32'h00000000;
assign filter_banks_24[13] = 32'h00000000;
assign filter_banks_24[14] = 32'h00000000;
assign filter_banks_24[15] = 32'h00000000;
assign filter_banks_24[16] = 32'h00000000;
assign filter_banks_24[17] = 32'h00000000;
assign filter_banks_24[18] = 32'h00000000;
assign filter_banks_24[19] = 32'h00000000;
assign filter_banks_24[20] = 32'h00000000;
assign filter_banks_24[21] = 32'h00000000;
assign filter_banks_24[22] = 32'h00000000;
assign filter_banks_24[23] = 32'h00000000;
assign filter_banks_24[24] = 32'h00000000;
assign filter_banks_24[25] = 32'h00000000;
assign filter_banks_24[26] = 32'h00000000;
assign filter_banks_24[27] = 32'h00000000;
assign filter_banks_24[28] = 32'h00000000;
assign filter_banks_24[29] = 32'h00000000;
assign filter_banks_24[30] = 32'h00000000;
assign filter_banks_24[31] = 32'h00000000;
assign filter_banks_24[32] = 32'h00000000;
assign filter_banks_24[33] = 32'h00000000;
assign filter_banks_24[34] = 32'h00000000;
assign filter_banks_24[35] = 32'h00000000;
assign filter_banks_24[36] = 32'h00000000;
assign filter_banks_24[37] = 32'h00000000;
assign filter_banks_24[38] = 32'h00000000;
assign filter_banks_24[39] = 32'h00000000;
assign filter_banks_24[40] = 32'h00000000;
assign filter_banks_24[41] = 32'h00000000;
assign filter_banks_24[42] = 32'h00000000;
assign filter_banks_24[43] = 32'h00000000;
assign filter_banks_24[44] = 32'h00000000;
assign filter_banks_24[45] = 32'h00000000;
assign filter_banks_24[46] = 32'h00000000;
assign filter_banks_24[47] = 32'h00000000;
assign filter_banks_24[48] = 32'h00000000;
assign filter_banks_24[49] = 32'h00000000;
assign filter_banks_24[50] = 32'h00000000;
assign filter_banks_24[51] = 32'h00000000;
assign filter_banks_24[52] = 32'h00000000;
assign filter_banks_24[53] = 32'h00000000;
assign filter_banks_24[54] = 32'h00000000;
assign filter_banks_24[55] = 32'h00000000;
assign filter_banks_24[56] = 32'h00000000;
assign filter_banks_24[57] = 32'h00000000;
assign filter_banks_24[58] = 32'h00000000;
assign filter_banks_24[59] = 32'h00000000;
assign filter_banks_24[60] = 32'h00000000;
assign filter_banks_24[61] = 32'h00000000;
assign filter_banks_24[62] = 32'h00000000;
assign filter_banks_24[63] = 32'h00000000;
assign filter_banks_24[64] = 32'h00000000;
assign filter_banks_24[65] = 32'h00000000;
assign filter_banks_24[66] = 32'h00000000;
assign filter_banks_24[67] = 32'h00000000;
assign filter_banks_24[68] = 32'h00000000;
assign filter_banks_24[69] = 32'h00000000;
assign filter_banks_24[70] = 32'h00000000;
assign filter_banks_24[71] = 32'h00000000;
assign filter_banks_24[72] = 32'h00000000;
assign filter_banks_24[73] = 32'h00000000;
assign filter_banks_24[74] = 32'h00000000;
assign filter_banks_24[75] = 32'h00000000;
assign filter_banks_24[76] = 32'h00000000;
assign filter_banks_24[77] = 32'h00000000;
assign filter_banks_24[78] = 32'h00000000;
assign filter_banks_24[79] = 32'h00000000;
assign filter_banks_24[80] = 32'h00000000;
assign filter_banks_24[81] = 32'h00000000;
assign filter_banks_24[82] = 32'h00000000;
assign filter_banks_24[83] = 32'h00000000;
assign filter_banks_24[84] = 32'h00000000;
assign filter_banks_24[85] = 32'h00000000;
assign filter_banks_24[86] = 32'h00000000;
assign filter_banks_24[87] = 32'h00000000;
assign filter_banks_24[88] = 32'h00000000;
assign filter_banks_24[89] = 32'h00000000;
assign filter_banks_24[90] = 32'h00000000;
assign filter_banks_24[91] = 32'h00000000;
assign filter_banks_24[92] = 32'h00000000;
assign filter_banks_24[93] = 32'h00000000;
assign filter_banks_24[94] = 32'h00000000;
assign filter_banks_24[95] = 32'h00000000;
assign filter_banks_24[96] = 32'h00000000;
assign filter_banks_24[97] = 32'h00000000;
assign filter_banks_24[98] = 32'h00000000;
assign filter_banks_24[99] = 32'h00000000;
assign filter_banks_24[100] = 32'h00000000;
assign filter_banks_24[101] = 32'h00000000;
assign filter_banks_24[102] = 32'h00000000;
assign filter_banks_24[103] = 32'h00000000;
assign filter_banks_24[104] = 32'h00000000;
assign filter_banks_24[105] = 32'h00000000;
assign filter_banks_24[106] = 32'h00000000;
assign filter_banks_24[107] = 32'h00000000;
assign filter_banks_24[108] = 32'h00000000;
assign filter_banks_24[109] = 32'h00000000;
assign filter_banks_24[110] = 32'h00000000;
assign filter_banks_24[111] = 32'h00000000;
assign filter_banks_24[112] = 32'h00000000;
assign filter_banks_24[113] = 32'h00000000;
assign filter_banks_24[114] = 32'h00000000;
assign filter_banks_24[115] = 32'h00000000;
assign filter_banks_24[116] = 32'h00000000;
assign filter_banks_24[117] = 32'h00000000;
assign filter_banks_24[118] = 32'h00000000;
assign filter_banks_24[119] = 32'h00000000;
assign filter_banks_24[120] = 32'h00000000;
assign filter_banks_24[121] = 32'h00000000;
assign filter_banks_24[122] = 32'h00000000;
assign filter_banks_24[123] = 32'h00000000;
assign filter_banks_24[124] = 32'h00000000;
assign filter_banks_24[125] = 32'h00000000;
assign filter_banks_24[126] = 32'h00000000;
assign filter_banks_24[127] = 32'h00000000;
assign filter_banks_24[128] = 32'h00000000;
assign filter_banks_24[129] = 32'h00000000;
assign filter_banks_24[130] = 32'h00000000;
assign filter_banks_24[131] = 32'h00000000;
assign filter_banks_24[132] = 32'h00000000;
assign filter_banks_24[133] = 32'h00000000;
assign filter_banks_24[134] = 32'h00000000;
assign filter_banks_24[135] = 32'h00000000;
assign filter_banks_24[136] = 32'h00000000;
assign filter_banks_24[137] = 32'h00000000;
assign filter_banks_24[138] = 32'h00000000;
assign filter_banks_24[139] = 32'h00000000;
assign filter_banks_24[140] = 32'h00000000;
assign filter_banks_24[141] = 32'h00000000;
assign filter_banks_24[142] = 32'h00000000;
assign filter_banks_24[143] = 32'h00000000;
assign filter_banks_24[144] = 32'h00000000;
assign filter_banks_24[145] = 32'h00000000;
assign filter_banks_24[146] = 32'h00000000;
assign filter_banks_24[147] = 32'h00000000;
assign filter_banks_24[148] = 32'h00000000;
assign filter_banks_24[149] = 32'h00000000;
assign filter_banks_24[150] = 32'h00000000;
assign filter_banks_24[151] = 32'h00000000;
assign filter_banks_24[152] = 32'h00000000;
assign filter_banks_24[153] = 32'h00000000;
assign filter_banks_24[154] = 32'h00000000;
assign filter_banks_24[155] = 32'h00000000;
assign filter_banks_24[156] = 32'h00000000;
assign filter_banks_24[157] = 32'h00000000;
assign filter_banks_24[158] = 32'h00000000;
assign filter_banks_24[159] = 32'h00000000;
assign filter_banks_24[160] = 32'h00000000;
assign filter_banks_24[161] = 32'h00000000;
assign filter_banks_24[162] = 32'h00000000;
assign filter_banks_24[163] = 32'h00000000;
assign filter_banks_24[164] = 32'h00000000;
assign filter_banks_24[165] = 32'h00000000;
assign filter_banks_24[166] = 32'h00000000;
assign filter_banks_24[167] = 32'h00000000;
assign filter_banks_24[168] = 32'h00000000;
assign filter_banks_24[169] = 32'h00000000;
assign filter_banks_24[170] = 32'h3d579436;
assign filter_banks_24[171] = 32'h3dd79436;
assign filter_banks_24[172] = 32'h3e21af28;
assign filter_banks_24[173] = 32'h3e579436;
assign filter_banks_24[174] = 32'h3e86bca2;
assign filter_banks_24[175] = 32'h3ea1af28;
assign filter_banks_24[176] = 32'h3ebca1af;
assign filter_banks_24[177] = 32'h3ed79436;
assign filter_banks_24[178] = 32'h3ef286bd;
assign filter_banks_24[179] = 32'h3f06bca2;
assign filter_banks_24[180] = 32'h3f1435e5;
assign filter_banks_24[181] = 32'h3f21af28;
assign filter_banks_24[182] = 32'h3f2f286c;
assign filter_banks_24[183] = 32'h3f3ca1af;
assign filter_banks_24[184] = 32'h3f4a1af3;
assign filter_banks_24[185] = 32'h3f579436;
assign filter_banks_24[186] = 32'h3f650d79;
assign filter_banks_24[187] = 32'h3f7286bd;
assign filter_banks_24[188] = 32'h3f800000;
assign filter_banks_24[189] = 32'h3f73cf3d;
assign filter_banks_24[190] = 32'h3f679e7a;
assign filter_banks_24[191] = 32'h3f5b6db7;
assign filter_banks_24[192] = 32'h3f4f3cf4;
assign filter_banks_24[193] = 32'h3f430c31;
assign filter_banks_24[194] = 32'h3f36db6e;
assign filter_banks_24[195] = 32'h3f2aaaab;
assign filter_banks_24[196] = 32'h3f1e79e8;
assign filter_banks_24[197] = 32'h3f124925;
assign filter_banks_24[198] = 32'h3f061862;
assign filter_banks_24[199] = 32'h3ef3cf3d;
assign filter_banks_24[200] = 32'h3edb6db7;
assign filter_banks_24[201] = 32'h3ec30c31;
assign filter_banks_24[202] = 32'h3eaaaaab;
assign filter_banks_24[203] = 32'h3e924925;
assign filter_banks_24[204] = 32'h3e73cf3d;
assign filter_banks_24[205] = 32'h3e430c31;
assign filter_banks_24[206] = 32'h3e124925;
assign filter_banks_24[207] = 32'h3dc30c31;
assign filter_banks_24[208] = 32'h3d430c31;
assign filter_banks_24[209] = 32'h00000000;
assign filter_banks_24[210] = 32'h00000000;
assign filter_banks_24[211] = 32'h00000000;
assign filter_banks_24[212] = 32'h00000000;
assign filter_banks_24[213] = 32'h00000000;
assign filter_banks_24[214] = 32'h00000000;
assign filter_banks_24[215] = 32'h00000000;
assign filter_banks_24[216] = 32'h00000000;
assign filter_banks_24[217] = 32'h00000000;
assign filter_banks_24[218] = 32'h00000000;
assign filter_banks_24[219] = 32'h00000000;
assign filter_banks_24[220] = 32'h00000000;
assign filter_banks_24[221] = 32'h00000000;
assign filter_banks_24[222] = 32'h00000000;
assign filter_banks_24[223] = 32'h00000000;
assign filter_banks_24[224] = 32'h00000000;
assign filter_banks_24[225] = 32'h00000000;
assign filter_banks_24[226] = 32'h00000000;
assign filter_banks_24[227] = 32'h00000000;
assign filter_banks_24[228] = 32'h00000000;
assign filter_banks_24[229] = 32'h00000000;
assign filter_banks_24[230] = 32'h00000000;
assign filter_banks_24[231] = 32'h00000000;
assign filter_banks_24[232] = 32'h00000000;
assign filter_banks_24[233] = 32'h00000000;
assign filter_banks_24[234] = 32'h00000000;
assign filter_banks_24[235] = 32'h00000000;
assign filter_banks_24[236] = 32'h00000000;
assign filter_banks_24[237] = 32'h00000000;
assign filter_banks_24[238] = 32'h00000000;
assign filter_banks_24[239] = 32'h00000000;
assign filter_banks_24[240] = 32'h00000000;
assign filter_banks_24[241] = 32'h00000000;
assign filter_banks_24[242] = 32'h00000000;
assign filter_banks_24[243] = 32'h00000000;
assign filter_banks_24[244] = 32'h00000000;
assign filter_banks_24[245] = 32'h00000000;
assign filter_banks_24[246] = 32'h00000000;
assign filter_banks_24[247] = 32'h00000000;
assign filter_banks_24[248] = 32'h00000000;
assign filter_banks_24[249] = 32'h00000000;
assign filter_banks_24[250] = 32'h00000000;
assign filter_banks_24[251] = 32'h00000000;
assign filter_banks_24[252] = 32'h00000000;
assign filter_banks_24[253] = 32'h00000000;
assign filter_banks_24[254] = 32'h00000000;
assign filter_banks_24[255] = 32'h00000000;
assign filter_banks_24[256] = 32'h00000000;
assign filter_banks_25[0] = 32'h00000000;
assign filter_banks_25[1] = 32'h00000000;
assign filter_banks_25[2] = 32'h00000000;
assign filter_banks_25[3] = 32'h00000000;
assign filter_banks_25[4] = 32'h00000000;
assign filter_banks_25[5] = 32'h00000000;
assign filter_banks_25[6] = 32'h00000000;
assign filter_banks_25[7] = 32'h00000000;
assign filter_banks_25[8] = 32'h00000000;
assign filter_banks_25[9] = 32'h00000000;
assign filter_banks_25[10] = 32'h00000000;
assign filter_banks_25[11] = 32'h00000000;
assign filter_banks_25[12] = 32'h00000000;
assign filter_banks_25[13] = 32'h00000000;
assign filter_banks_25[14] = 32'h00000000;
assign filter_banks_25[15] = 32'h00000000;
assign filter_banks_25[16] = 32'h00000000;
assign filter_banks_25[17] = 32'h00000000;
assign filter_banks_25[18] = 32'h00000000;
assign filter_banks_25[19] = 32'h00000000;
assign filter_banks_25[20] = 32'h00000000;
assign filter_banks_25[21] = 32'h00000000;
assign filter_banks_25[22] = 32'h00000000;
assign filter_banks_25[23] = 32'h00000000;
assign filter_banks_25[24] = 32'h00000000;
assign filter_banks_25[25] = 32'h00000000;
assign filter_banks_25[26] = 32'h00000000;
assign filter_banks_25[27] = 32'h00000000;
assign filter_banks_25[28] = 32'h00000000;
assign filter_banks_25[29] = 32'h00000000;
assign filter_banks_25[30] = 32'h00000000;
assign filter_banks_25[31] = 32'h00000000;
assign filter_banks_25[32] = 32'h00000000;
assign filter_banks_25[33] = 32'h00000000;
assign filter_banks_25[34] = 32'h00000000;
assign filter_banks_25[35] = 32'h00000000;
assign filter_banks_25[36] = 32'h00000000;
assign filter_banks_25[37] = 32'h00000000;
assign filter_banks_25[38] = 32'h00000000;
assign filter_banks_25[39] = 32'h00000000;
assign filter_banks_25[40] = 32'h00000000;
assign filter_banks_25[41] = 32'h00000000;
assign filter_banks_25[42] = 32'h00000000;
assign filter_banks_25[43] = 32'h00000000;
assign filter_banks_25[44] = 32'h00000000;
assign filter_banks_25[45] = 32'h00000000;
assign filter_banks_25[46] = 32'h00000000;
assign filter_banks_25[47] = 32'h00000000;
assign filter_banks_25[48] = 32'h00000000;
assign filter_banks_25[49] = 32'h00000000;
assign filter_banks_25[50] = 32'h00000000;
assign filter_banks_25[51] = 32'h00000000;
assign filter_banks_25[52] = 32'h00000000;
assign filter_banks_25[53] = 32'h00000000;
assign filter_banks_25[54] = 32'h00000000;
assign filter_banks_25[55] = 32'h00000000;
assign filter_banks_25[56] = 32'h00000000;
assign filter_banks_25[57] = 32'h00000000;
assign filter_banks_25[58] = 32'h00000000;
assign filter_banks_25[59] = 32'h00000000;
assign filter_banks_25[60] = 32'h00000000;
assign filter_banks_25[61] = 32'h00000000;
assign filter_banks_25[62] = 32'h00000000;
assign filter_banks_25[63] = 32'h00000000;
assign filter_banks_25[64] = 32'h00000000;
assign filter_banks_25[65] = 32'h00000000;
assign filter_banks_25[66] = 32'h00000000;
assign filter_banks_25[67] = 32'h00000000;
assign filter_banks_25[68] = 32'h00000000;
assign filter_banks_25[69] = 32'h00000000;
assign filter_banks_25[70] = 32'h00000000;
assign filter_banks_25[71] = 32'h00000000;
assign filter_banks_25[72] = 32'h00000000;
assign filter_banks_25[73] = 32'h00000000;
assign filter_banks_25[74] = 32'h00000000;
assign filter_banks_25[75] = 32'h00000000;
assign filter_banks_25[76] = 32'h00000000;
assign filter_banks_25[77] = 32'h00000000;
assign filter_banks_25[78] = 32'h00000000;
assign filter_banks_25[79] = 32'h00000000;
assign filter_banks_25[80] = 32'h00000000;
assign filter_banks_25[81] = 32'h00000000;
assign filter_banks_25[82] = 32'h00000000;
assign filter_banks_25[83] = 32'h00000000;
assign filter_banks_25[84] = 32'h00000000;
assign filter_banks_25[85] = 32'h00000000;
assign filter_banks_25[86] = 32'h00000000;
assign filter_banks_25[87] = 32'h00000000;
assign filter_banks_25[88] = 32'h00000000;
assign filter_banks_25[89] = 32'h00000000;
assign filter_banks_25[90] = 32'h00000000;
assign filter_banks_25[91] = 32'h00000000;
assign filter_banks_25[92] = 32'h00000000;
assign filter_banks_25[93] = 32'h00000000;
assign filter_banks_25[94] = 32'h00000000;
assign filter_banks_25[95] = 32'h00000000;
assign filter_banks_25[96] = 32'h00000000;
assign filter_banks_25[97] = 32'h00000000;
assign filter_banks_25[98] = 32'h00000000;
assign filter_banks_25[99] = 32'h00000000;
assign filter_banks_25[100] = 32'h00000000;
assign filter_banks_25[101] = 32'h00000000;
assign filter_banks_25[102] = 32'h00000000;
assign filter_banks_25[103] = 32'h00000000;
assign filter_banks_25[104] = 32'h00000000;
assign filter_banks_25[105] = 32'h00000000;
assign filter_banks_25[106] = 32'h00000000;
assign filter_banks_25[107] = 32'h00000000;
assign filter_banks_25[108] = 32'h00000000;
assign filter_banks_25[109] = 32'h00000000;
assign filter_banks_25[110] = 32'h00000000;
assign filter_banks_25[111] = 32'h00000000;
assign filter_banks_25[112] = 32'h00000000;
assign filter_banks_25[113] = 32'h00000000;
assign filter_banks_25[114] = 32'h00000000;
assign filter_banks_25[115] = 32'h00000000;
assign filter_banks_25[116] = 32'h00000000;
assign filter_banks_25[117] = 32'h00000000;
assign filter_banks_25[118] = 32'h00000000;
assign filter_banks_25[119] = 32'h00000000;
assign filter_banks_25[120] = 32'h00000000;
assign filter_banks_25[121] = 32'h00000000;
assign filter_banks_25[122] = 32'h00000000;
assign filter_banks_25[123] = 32'h00000000;
assign filter_banks_25[124] = 32'h00000000;
assign filter_banks_25[125] = 32'h00000000;
assign filter_banks_25[126] = 32'h00000000;
assign filter_banks_25[127] = 32'h00000000;
assign filter_banks_25[128] = 32'h00000000;
assign filter_banks_25[129] = 32'h00000000;
assign filter_banks_25[130] = 32'h00000000;
assign filter_banks_25[131] = 32'h00000000;
assign filter_banks_25[132] = 32'h00000000;
assign filter_banks_25[133] = 32'h00000000;
assign filter_banks_25[134] = 32'h00000000;
assign filter_banks_25[135] = 32'h00000000;
assign filter_banks_25[136] = 32'h00000000;
assign filter_banks_25[137] = 32'h00000000;
assign filter_banks_25[138] = 32'h00000000;
assign filter_banks_25[139] = 32'h00000000;
assign filter_banks_25[140] = 32'h00000000;
assign filter_banks_25[141] = 32'h00000000;
assign filter_banks_25[142] = 32'h00000000;
assign filter_banks_25[143] = 32'h00000000;
assign filter_banks_25[144] = 32'h00000000;
assign filter_banks_25[145] = 32'h00000000;
assign filter_banks_25[146] = 32'h00000000;
assign filter_banks_25[147] = 32'h00000000;
assign filter_banks_25[148] = 32'h00000000;
assign filter_banks_25[149] = 32'h00000000;
assign filter_banks_25[150] = 32'h00000000;
assign filter_banks_25[151] = 32'h00000000;
assign filter_banks_25[152] = 32'h00000000;
assign filter_banks_25[153] = 32'h00000000;
assign filter_banks_25[154] = 32'h00000000;
assign filter_banks_25[155] = 32'h00000000;
assign filter_banks_25[156] = 32'h00000000;
assign filter_banks_25[157] = 32'h00000000;
assign filter_banks_25[158] = 32'h00000000;
assign filter_banks_25[159] = 32'h00000000;
assign filter_banks_25[160] = 32'h00000000;
assign filter_banks_25[161] = 32'h00000000;
assign filter_banks_25[162] = 32'h00000000;
assign filter_banks_25[163] = 32'h00000000;
assign filter_banks_25[164] = 32'h00000000;
assign filter_banks_25[165] = 32'h00000000;
assign filter_banks_25[166] = 32'h00000000;
assign filter_banks_25[167] = 32'h00000000;
assign filter_banks_25[168] = 32'h00000000;
assign filter_banks_25[169] = 32'h00000000;
assign filter_banks_25[170] = 32'h00000000;
assign filter_banks_25[171] = 32'h00000000;
assign filter_banks_25[172] = 32'h00000000;
assign filter_banks_25[173] = 32'h00000000;
assign filter_banks_25[174] = 32'h00000000;
assign filter_banks_25[175] = 32'h00000000;
assign filter_banks_25[176] = 32'h00000000;
assign filter_banks_25[177] = 32'h00000000;
assign filter_banks_25[178] = 32'h00000000;
assign filter_banks_25[179] = 32'h00000000;
assign filter_banks_25[180] = 32'h00000000;
assign filter_banks_25[181] = 32'h00000000;
assign filter_banks_25[182] = 32'h00000000;
assign filter_banks_25[183] = 32'h00000000;
assign filter_banks_25[184] = 32'h00000000;
assign filter_banks_25[185] = 32'h00000000;
assign filter_banks_25[186] = 32'h00000000;
assign filter_banks_25[187] = 32'h00000000;
assign filter_banks_25[188] = 32'h00000000;
assign filter_banks_25[189] = 32'h3d430c31;
assign filter_banks_25[190] = 32'h3dc30c31;
assign filter_banks_25[191] = 32'h3e124925;
assign filter_banks_25[192] = 32'h3e430c31;
assign filter_banks_25[193] = 32'h3e73cf3d;
assign filter_banks_25[194] = 32'h3e924925;
assign filter_banks_25[195] = 32'h3eaaaaab;
assign filter_banks_25[196] = 32'h3ec30c31;
assign filter_banks_25[197] = 32'h3edb6db7;
assign filter_banks_25[198] = 32'h3ef3cf3d;
assign filter_banks_25[199] = 32'h3f061862;
assign filter_banks_25[200] = 32'h3f124925;
assign filter_banks_25[201] = 32'h3f1e79e8;
assign filter_banks_25[202] = 32'h3f2aaaab;
assign filter_banks_25[203] = 32'h3f36db6e;
assign filter_banks_25[204] = 32'h3f430c31;
assign filter_banks_25[205] = 32'h3f4f3cf4;
assign filter_banks_25[206] = 32'h3f5b6db7;
assign filter_banks_25[207] = 32'h3f679e7a;
assign filter_banks_25[208] = 32'h3f73cf3d;
assign filter_banks_25[209] = 32'h3f800000;
assign filter_banks_25[210] = 32'h3f745d17;
assign filter_banks_25[211] = 32'h3f68ba2f;
assign filter_banks_25[212] = 32'h3f5d1746;
assign filter_banks_25[213] = 32'h3f51745d;
assign filter_banks_25[214] = 32'h3f45d174;
assign filter_banks_25[215] = 32'h3f3a2e8c;
assign filter_banks_25[216] = 32'h3f2e8ba3;
assign filter_banks_25[217] = 32'h3f22e8ba;
assign filter_banks_25[218] = 32'h3f1745d1;
assign filter_banks_25[219] = 32'h3f0ba2e9;
assign filter_banks_25[220] = 32'h3f000000;
assign filter_banks_25[221] = 32'h3ee8ba2f;
assign filter_banks_25[222] = 32'h3ed1745d;
assign filter_banks_25[223] = 32'h3eba2e8c;
assign filter_banks_25[224] = 32'h3ea2e8ba;
assign filter_banks_25[225] = 32'h3e8ba2e9;
assign filter_banks_25[226] = 32'h3e68ba2f;
assign filter_banks_25[227] = 32'h3e3a2e8c;
assign filter_banks_25[228] = 32'h3e0ba2e9;
assign filter_banks_25[229] = 32'h3dba2e8c;
assign filter_banks_25[230] = 32'h3d3a2e8c;
assign filter_banks_25[231] = 32'h00000000;
assign filter_banks_25[232] = 32'h00000000;
assign filter_banks_25[233] = 32'h00000000;
assign filter_banks_25[234] = 32'h00000000;
assign filter_banks_25[235] = 32'h00000000;
assign filter_banks_25[236] = 32'h00000000;
assign filter_banks_25[237] = 32'h00000000;
assign filter_banks_25[238] = 32'h00000000;
assign filter_banks_25[239] = 32'h00000000;
assign filter_banks_25[240] = 32'h00000000;
assign filter_banks_25[241] = 32'h00000000;
assign filter_banks_25[242] = 32'h00000000;
assign filter_banks_25[243] = 32'h00000000;
assign filter_banks_25[244] = 32'h00000000;
assign filter_banks_25[245] = 32'h00000000;
assign filter_banks_25[246] = 32'h00000000;
assign filter_banks_25[247] = 32'h00000000;
assign filter_banks_25[248] = 32'h00000000;
assign filter_banks_25[249] = 32'h00000000;
assign filter_banks_25[250] = 32'h00000000;
assign filter_banks_25[251] = 32'h00000000;
assign filter_banks_25[252] = 32'h00000000;
assign filter_banks_25[253] = 32'h00000000;
assign filter_banks_25[254] = 32'h00000000;
assign filter_banks_25[255] = 32'h00000000;
assign filter_banks_25[256] = 32'h00000000;
assign filter_banks_26[0] = 32'h00000000;
assign filter_banks_26[1] = 32'h00000000;
assign filter_banks_26[2] = 32'h00000000;
assign filter_banks_26[3] = 32'h00000000;
assign filter_banks_26[4] = 32'h00000000;
assign filter_banks_26[5] = 32'h00000000;
assign filter_banks_26[6] = 32'h00000000;
assign filter_banks_26[7] = 32'h00000000;
assign filter_banks_26[8] = 32'h00000000;
assign filter_banks_26[9] = 32'h00000000;
assign filter_banks_26[10] = 32'h00000000;
assign filter_banks_26[11] = 32'h00000000;
assign filter_banks_26[12] = 32'h00000000;
assign filter_banks_26[13] = 32'h00000000;
assign filter_banks_26[14] = 32'h00000000;
assign filter_banks_26[15] = 32'h00000000;
assign filter_banks_26[16] = 32'h00000000;
assign filter_banks_26[17] = 32'h00000000;
assign filter_banks_26[18] = 32'h00000000;
assign filter_banks_26[19] = 32'h00000000;
assign filter_banks_26[20] = 32'h00000000;
assign filter_banks_26[21] = 32'h00000000;
assign filter_banks_26[22] = 32'h00000000;
assign filter_banks_26[23] = 32'h00000000;
assign filter_banks_26[24] = 32'h00000000;
assign filter_banks_26[25] = 32'h00000000;
assign filter_banks_26[26] = 32'h00000000;
assign filter_banks_26[27] = 32'h00000000;
assign filter_banks_26[28] = 32'h00000000;
assign filter_banks_26[29] = 32'h00000000;
assign filter_banks_26[30] = 32'h00000000;
assign filter_banks_26[31] = 32'h00000000;
assign filter_banks_26[32] = 32'h00000000;
assign filter_banks_26[33] = 32'h00000000;
assign filter_banks_26[34] = 32'h00000000;
assign filter_banks_26[35] = 32'h00000000;
assign filter_banks_26[36] = 32'h00000000;
assign filter_banks_26[37] = 32'h00000000;
assign filter_banks_26[38] = 32'h00000000;
assign filter_banks_26[39] = 32'h00000000;
assign filter_banks_26[40] = 32'h00000000;
assign filter_banks_26[41] = 32'h00000000;
assign filter_banks_26[42] = 32'h00000000;
assign filter_banks_26[43] = 32'h00000000;
assign filter_banks_26[44] = 32'h00000000;
assign filter_banks_26[45] = 32'h00000000;
assign filter_banks_26[46] = 32'h00000000;
assign filter_banks_26[47] = 32'h00000000;
assign filter_banks_26[48] = 32'h00000000;
assign filter_banks_26[49] = 32'h00000000;
assign filter_banks_26[50] = 32'h00000000;
assign filter_banks_26[51] = 32'h00000000;
assign filter_banks_26[52] = 32'h00000000;
assign filter_banks_26[53] = 32'h00000000;
assign filter_banks_26[54] = 32'h00000000;
assign filter_banks_26[55] = 32'h00000000;
assign filter_banks_26[56] = 32'h00000000;
assign filter_banks_26[57] = 32'h00000000;
assign filter_banks_26[58] = 32'h00000000;
assign filter_banks_26[59] = 32'h00000000;
assign filter_banks_26[60] = 32'h00000000;
assign filter_banks_26[61] = 32'h00000000;
assign filter_banks_26[62] = 32'h00000000;
assign filter_banks_26[63] = 32'h00000000;
assign filter_banks_26[64] = 32'h00000000;
assign filter_banks_26[65] = 32'h00000000;
assign filter_banks_26[66] = 32'h00000000;
assign filter_banks_26[67] = 32'h00000000;
assign filter_banks_26[68] = 32'h00000000;
assign filter_banks_26[69] = 32'h00000000;
assign filter_banks_26[70] = 32'h00000000;
assign filter_banks_26[71] = 32'h00000000;
assign filter_banks_26[72] = 32'h00000000;
assign filter_banks_26[73] = 32'h00000000;
assign filter_banks_26[74] = 32'h00000000;
assign filter_banks_26[75] = 32'h00000000;
assign filter_banks_26[76] = 32'h00000000;
assign filter_banks_26[77] = 32'h00000000;
assign filter_banks_26[78] = 32'h00000000;
assign filter_banks_26[79] = 32'h00000000;
assign filter_banks_26[80] = 32'h00000000;
assign filter_banks_26[81] = 32'h00000000;
assign filter_banks_26[82] = 32'h00000000;
assign filter_banks_26[83] = 32'h00000000;
assign filter_banks_26[84] = 32'h00000000;
assign filter_banks_26[85] = 32'h00000000;
assign filter_banks_26[86] = 32'h00000000;
assign filter_banks_26[87] = 32'h00000000;
assign filter_banks_26[88] = 32'h00000000;
assign filter_banks_26[89] = 32'h00000000;
assign filter_banks_26[90] = 32'h00000000;
assign filter_banks_26[91] = 32'h00000000;
assign filter_banks_26[92] = 32'h00000000;
assign filter_banks_26[93] = 32'h00000000;
assign filter_banks_26[94] = 32'h00000000;
assign filter_banks_26[95] = 32'h00000000;
assign filter_banks_26[96] = 32'h00000000;
assign filter_banks_26[97] = 32'h00000000;
assign filter_banks_26[98] = 32'h00000000;
assign filter_banks_26[99] = 32'h00000000;
assign filter_banks_26[100] = 32'h00000000;
assign filter_banks_26[101] = 32'h00000000;
assign filter_banks_26[102] = 32'h00000000;
assign filter_banks_26[103] = 32'h00000000;
assign filter_banks_26[104] = 32'h00000000;
assign filter_banks_26[105] = 32'h00000000;
assign filter_banks_26[106] = 32'h00000000;
assign filter_banks_26[107] = 32'h00000000;
assign filter_banks_26[108] = 32'h00000000;
assign filter_banks_26[109] = 32'h00000000;
assign filter_banks_26[110] = 32'h00000000;
assign filter_banks_26[111] = 32'h00000000;
assign filter_banks_26[112] = 32'h00000000;
assign filter_banks_26[113] = 32'h00000000;
assign filter_banks_26[114] = 32'h00000000;
assign filter_banks_26[115] = 32'h00000000;
assign filter_banks_26[116] = 32'h00000000;
assign filter_banks_26[117] = 32'h00000000;
assign filter_banks_26[118] = 32'h00000000;
assign filter_banks_26[119] = 32'h00000000;
assign filter_banks_26[120] = 32'h00000000;
assign filter_banks_26[121] = 32'h00000000;
assign filter_banks_26[122] = 32'h00000000;
assign filter_banks_26[123] = 32'h00000000;
assign filter_banks_26[124] = 32'h00000000;
assign filter_banks_26[125] = 32'h00000000;
assign filter_banks_26[126] = 32'h00000000;
assign filter_banks_26[127] = 32'h00000000;
assign filter_banks_26[128] = 32'h00000000;
assign filter_banks_26[129] = 32'h00000000;
assign filter_banks_26[130] = 32'h00000000;
assign filter_banks_26[131] = 32'h00000000;
assign filter_banks_26[132] = 32'h00000000;
assign filter_banks_26[133] = 32'h00000000;
assign filter_banks_26[134] = 32'h00000000;
assign filter_banks_26[135] = 32'h00000000;
assign filter_banks_26[136] = 32'h00000000;
assign filter_banks_26[137] = 32'h00000000;
assign filter_banks_26[138] = 32'h00000000;
assign filter_banks_26[139] = 32'h00000000;
assign filter_banks_26[140] = 32'h00000000;
assign filter_banks_26[141] = 32'h00000000;
assign filter_banks_26[142] = 32'h00000000;
assign filter_banks_26[143] = 32'h00000000;
assign filter_banks_26[144] = 32'h00000000;
assign filter_banks_26[145] = 32'h00000000;
assign filter_banks_26[146] = 32'h00000000;
assign filter_banks_26[147] = 32'h00000000;
assign filter_banks_26[148] = 32'h00000000;
assign filter_banks_26[149] = 32'h00000000;
assign filter_banks_26[150] = 32'h00000000;
assign filter_banks_26[151] = 32'h00000000;
assign filter_banks_26[152] = 32'h00000000;
assign filter_banks_26[153] = 32'h00000000;
assign filter_banks_26[154] = 32'h00000000;
assign filter_banks_26[155] = 32'h00000000;
assign filter_banks_26[156] = 32'h00000000;
assign filter_banks_26[157] = 32'h00000000;
assign filter_banks_26[158] = 32'h00000000;
assign filter_banks_26[159] = 32'h00000000;
assign filter_banks_26[160] = 32'h00000000;
assign filter_banks_26[161] = 32'h00000000;
assign filter_banks_26[162] = 32'h00000000;
assign filter_banks_26[163] = 32'h00000000;
assign filter_banks_26[164] = 32'h00000000;
assign filter_banks_26[165] = 32'h00000000;
assign filter_banks_26[166] = 32'h00000000;
assign filter_banks_26[167] = 32'h00000000;
assign filter_banks_26[168] = 32'h00000000;
assign filter_banks_26[169] = 32'h00000000;
assign filter_banks_26[170] = 32'h00000000;
assign filter_banks_26[171] = 32'h00000000;
assign filter_banks_26[172] = 32'h00000000;
assign filter_banks_26[173] = 32'h00000000;
assign filter_banks_26[174] = 32'h00000000;
assign filter_banks_26[175] = 32'h00000000;
assign filter_banks_26[176] = 32'h00000000;
assign filter_banks_26[177] = 32'h00000000;
assign filter_banks_26[178] = 32'h00000000;
assign filter_banks_26[179] = 32'h00000000;
assign filter_banks_26[180] = 32'h00000000;
assign filter_banks_26[181] = 32'h00000000;
assign filter_banks_26[182] = 32'h00000000;
assign filter_banks_26[183] = 32'h00000000;
assign filter_banks_26[184] = 32'h00000000;
assign filter_banks_26[185] = 32'h00000000;
assign filter_banks_26[186] = 32'h00000000;
assign filter_banks_26[187] = 32'h00000000;
assign filter_banks_26[188] = 32'h00000000;
assign filter_banks_26[189] = 32'h00000000;
assign filter_banks_26[190] = 32'h00000000;
assign filter_banks_26[191] = 32'h00000000;
assign filter_banks_26[192] = 32'h00000000;
assign filter_banks_26[193] = 32'h00000000;
assign filter_banks_26[194] = 32'h00000000;
assign filter_banks_26[195] = 32'h00000000;
assign filter_banks_26[196] = 32'h00000000;
assign filter_banks_26[197] = 32'h00000000;
assign filter_banks_26[198] = 32'h00000000;
assign filter_banks_26[199] = 32'h00000000;
assign filter_banks_26[200] = 32'h00000000;
assign filter_banks_26[201] = 32'h00000000;
assign filter_banks_26[202] = 32'h00000000;
assign filter_banks_26[203] = 32'h00000000;
assign filter_banks_26[204] = 32'h00000000;
assign filter_banks_26[205] = 32'h00000000;
assign filter_banks_26[206] = 32'h00000000;
assign filter_banks_26[207] = 32'h00000000;
assign filter_banks_26[208] = 32'h00000000;
assign filter_banks_26[209] = 32'h00000000;
assign filter_banks_26[210] = 32'h3d3a2e8c;
assign filter_banks_26[211] = 32'h3dba2e8c;
assign filter_banks_26[212] = 32'h3e0ba2e9;
assign filter_banks_26[213] = 32'h3e3a2e8c;
assign filter_banks_26[214] = 32'h3e68ba2f;
assign filter_banks_26[215] = 32'h3e8ba2e9;
assign filter_banks_26[216] = 32'h3ea2e8ba;
assign filter_banks_26[217] = 32'h3eba2e8c;
assign filter_banks_26[218] = 32'h3ed1745d;
assign filter_banks_26[219] = 32'h3ee8ba2f;
assign filter_banks_26[220] = 32'h3f000000;
assign filter_banks_26[221] = 32'h3f0ba2e9;
assign filter_banks_26[222] = 32'h3f1745d1;
assign filter_banks_26[223] = 32'h3f22e8ba;
assign filter_banks_26[224] = 32'h3f2e8ba3;
assign filter_banks_26[225] = 32'h3f3a2e8c;
assign filter_banks_26[226] = 32'h3f45d174;
assign filter_banks_26[227] = 32'h3f51745d;
assign filter_banks_26[228] = 32'h3f5d1746;
assign filter_banks_26[229] = 32'h3f68ba2f;
assign filter_banks_26[230] = 32'h3f745d17;
assign filter_banks_26[231] = 32'h3f800000;
assign filter_banks_26[232] = 32'h3f75c28f;
assign filter_banks_26[233] = 32'h3f6b851f;
assign filter_banks_26[234] = 32'h3f6147ae;
assign filter_banks_26[235] = 32'h3f570a3d;
assign filter_banks_26[236] = 32'h3f4ccccd;
assign filter_banks_26[237] = 32'h3f428f5c;
assign filter_banks_26[238] = 32'h3f3851ec;
assign filter_banks_26[239] = 32'h3f2e147b;
assign filter_banks_26[240] = 32'h3f23d70a;
assign filter_banks_26[241] = 32'h3f19999a;
assign filter_banks_26[242] = 32'h3f0f5c29;
assign filter_banks_26[243] = 32'h3f051eb8;
assign filter_banks_26[244] = 32'h3ef5c28f;
assign filter_banks_26[245] = 32'h3ee147ae;
assign filter_banks_26[246] = 32'h3ecccccd;
assign filter_banks_26[247] = 32'h3eb851ec;
assign filter_banks_26[248] = 32'h3ea3d70a;
assign filter_banks_26[249] = 32'h3e8f5c29;
assign filter_banks_26[250] = 32'h3e75c28f;
assign filter_banks_26[251] = 32'h3e4ccccd;
assign filter_banks_26[252] = 32'h3e23d70a;
assign filter_banks_26[253] = 32'h3df5c28f;
assign filter_banks_26[254] = 32'h3da3d70a;
assign filter_banks_26[255] = 32'h3d23d70a;
assign filter_banks_26[256] = 32'h00000000;

    floating_point_mult_non_blocking m1_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[0]),
        .s_axis_b_tdata(reg_fb_1),
        .m_axis_result_tvalid(tvalid_res_mult_fb[0]),
        .m_axis_result_tdata(res_mult_fb_1)
    );
    
    floating_point_mult_non_blocking m2_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[1]),
        .s_axis_b_tdata(reg_fb_2),
        .m_axis_result_tvalid(tvalid_res_mult_fb[1]),
        .m_axis_result_tdata(res_mult_fb_2)
    );
    
    floating_point_mult_non_blocking m3_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[2]),
        .s_axis_b_tdata(reg_fb_3),
        .m_axis_result_tvalid(tvalid_res_mult_fb[2]),
        .m_axis_result_tdata(res_mult_fb_3)
    );
    
    floating_point_mult_non_blocking m4_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[3]),
        .s_axis_b_tdata(reg_fb_4),
        .m_axis_result_tvalid(tvalid_res_mult_fb[3]),
        .m_axis_result_tdata(res_mult_fb_4)
    );
    
    floating_point_mult_non_blocking m5_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[4]),
        .s_axis_b_tdata(reg_fb_5),
        .m_axis_result_tvalid(tvalid_res_mult_fb[4]),
        .m_axis_result_tdata(res_mult_fb_5)
    );
    
    floating_point_mult_non_blocking m6_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[5]),
        .s_axis_b_tdata(reg_fb_6),
        .m_axis_result_tvalid(tvalid_res_mult_fb[5]),
        .m_axis_result_tdata(res_mult_fb_6)
    );
    
    floating_point_mult_non_blocking m7_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[6]),
        .s_axis_b_tdata(reg_fb_7),
        .m_axis_result_tvalid(tvalid_res_mult_fb[6]),
        .m_axis_result_tdata(res_mult_fb_7)
    );
    
    floating_point_mult_non_blocking m8_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[7]),
        .s_axis_b_tdata(reg_fb_8),
        .m_axis_result_tvalid(tvalid_res_mult_fb[7]),
        .m_axis_result_tdata(res_mult_fb_8)
    );
    
    floating_point_mult_non_blocking m9_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[8]),
        .s_axis_b_tdata(reg_fb_9),
        .m_axis_result_tvalid(tvalid_res_mult_fb[8]),
        .m_axis_result_tdata(res_mult_fb_9)
    );
    
    floating_point_mult_non_blocking m10_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[9]),
        .s_axis_b_tdata(reg_fb_10),
        .m_axis_result_tvalid(tvalid_res_mult_fb[9]),
        .m_axis_result_tdata(res_mult_fb_10)
    );
    
    floating_point_mult_non_blocking m11_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[10]),
        .s_axis_b_tdata(reg_fb_11),
        .m_axis_result_tvalid(tvalid_res_mult_fb[10]),
        .m_axis_result_tdata(res_mult_fb_11)
    );
    
    floating_point_mult_non_blocking m12_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[11]),
        .s_axis_b_tdata(reg_fb_12),
        .m_axis_result_tvalid(tvalid_res_mult_fb[11]),
        .m_axis_result_tdata(res_mult_fb_12)
    );
    
    floating_point_mult_non_blocking m13_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[12]),
        .s_axis_b_tdata(reg_fb_13),
        .m_axis_result_tvalid(tvalid_res_mult_fb[12]),
        .m_axis_result_tdata(res_mult_fb_13)
    );
    
    floating_point_mult_non_blocking m14_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[13]),
        .s_axis_b_tdata(reg_fb_14),
        .m_axis_result_tvalid(tvalid_res_mult_fb[13]),
        .m_axis_result_tdata(res_mult_fb_14)
    );
    
    floating_point_mult_non_blocking m15_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[14]),
        .s_axis_b_tdata(reg_fb_15),
        .m_axis_result_tvalid(tvalid_res_mult_fb[14]),
        .m_axis_result_tdata(res_mult_fb_15)
    );
    
    floating_point_mult_non_blocking m16_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[15]),
        .s_axis_b_tdata(reg_fb_16),
        .m_axis_result_tvalid(tvalid_res_mult_fb[15]),
        .m_axis_result_tdata(res_mult_fb_16)
    );
    
    floating_point_mult_non_blocking m17_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[16]),
        .s_axis_b_tdata(reg_fb_17),
        .m_axis_result_tvalid(tvalid_res_mult_fb[16]),
        .m_axis_result_tdata(res_mult_fb_17)
    );
    
    floating_point_mult_non_blocking m18_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[17]),
        .s_axis_b_tdata(reg_fb_18),
        .m_axis_result_tvalid(tvalid_res_mult_fb[17]),
        .m_axis_result_tdata(res_mult_fb_18)
    );
    
    floating_point_mult_non_blocking m19_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[18]),
        .s_axis_b_tdata(reg_fb_19),
        .m_axis_result_tvalid(tvalid_res_mult_fb[18]),
        .m_axis_result_tdata(res_mult_fb_19)
    );
    
    floating_point_mult_non_blocking m20_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[19]),
        .s_axis_b_tdata(reg_fb_20),
        .m_axis_result_tvalid(tvalid_res_mult_fb[19]),
        .m_axis_result_tdata(res_mult_fb_20)
    );
    
    floating_point_mult_non_blocking m21_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[20]),
        .s_axis_b_tdata(reg_fb_21),
        .m_axis_result_tvalid(tvalid_res_mult_fb[20]),
        .m_axis_result_tdata(res_mult_fb_21)
    );
    
    floating_point_mult_non_blocking m22_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[21]),
        .s_axis_b_tdata(reg_fb_22),
        .m_axis_result_tvalid(tvalid_res_mult_fb[21]),
        .m_axis_result_tdata(res_mult_fb_22)
    );
    
    floating_point_mult_non_blocking m23_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[22]),
        .s_axis_b_tdata(reg_fb_23),
        .m_axis_result_tvalid(tvalid_res_mult_fb[22]),
        .m_axis_result_tdata(res_mult_fb_23)
    );
    
    floating_point_mult_non_blocking m24_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[23]),
        .s_axis_b_tdata(reg_fb_24),
        .m_axis_result_tvalid(tvalid_res_mult_fb[23]),
        .m_axis_result_tdata(res_mult_fb_24)
    );
    
    floating_point_mult_non_blocking m25_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[24]),
        .s_axis_b_tdata(reg_fb_25),
        .m_axis_result_tvalid(tvalid_res_mult_fb[24]),
        .m_axis_result_tdata(res_mult_fb_25)
    );
    
    floating_point_mult_non_blocking m26_mult_fb (
        .s_axis_a_tvalid(tvalid_powspectr),
        .s_axis_a_tdata(powspectr_temp),
        .s_axis_b_tvalid(tvalid_reg_fb[25]),
        .s_axis_b_tdata(reg_fb_26),
        .m_axis_result_tvalid(tvalid_res_mult_fb[25]),
        .m_axis_result_tdata(res_mult_fb_26)
    );
    
    floating_point_add_non_blocking m1_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[0]),
        .s_axis_a_tdata(res_mult_fb_1),
        .s_axis_b_tvalid(tvalid_out_acc[0]),
        .s_axis_b_tdata(out_acc_1),
        .m_axis_result_tvalid(tvalid_res_add_fb[0]),
        .m_axis_result_tdata(res_add_fb_1)
    );
    
    floating_point_add_non_blocking m2_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[1]),
        .s_axis_a_tdata(res_mult_fb_2),
        .s_axis_b_tvalid(tvalid_out_acc[1]),
        .s_axis_b_tdata(out_acc_2),
        .m_axis_result_tvalid(tvalid_res_add_fb[1]),
        .m_axis_result_tdata(res_add_fb_2)
    );
    
    floating_point_add_non_blocking m3_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[2]),
        .s_axis_a_tdata(res_mult_fb_3),
        .s_axis_b_tvalid(tvalid_out_acc[2]),
        .s_axis_b_tdata(out_acc_3),
        .m_axis_result_tvalid(tvalid_res_add_fb[2]),
        .m_axis_result_tdata(res_add_fb_3)
    );
    
    floating_point_add_non_blocking m4_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[3]),
        .s_axis_a_tdata(res_mult_fb_4),
        .s_axis_b_tvalid(tvalid_out_acc[3]),
        .s_axis_b_tdata(out_acc_4),
        .m_axis_result_tvalid(tvalid_res_add_fb[3]),
        .m_axis_result_tdata(res_add_fb_4)
    );
    
    floating_point_add_non_blocking m5_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[4]),
        .s_axis_a_tdata(res_mult_fb_5),
        .s_axis_b_tvalid(tvalid_out_acc[4]),
        .s_axis_b_tdata(out_acc_5),
        .m_axis_result_tvalid(tvalid_res_add_fb[4]),
        .m_axis_result_tdata(res_add_fb_5)
    );
    
    floating_point_add_non_blocking m6_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[5]),
        .s_axis_a_tdata(res_mult_fb_6),
        .s_axis_b_tvalid(tvalid_out_acc[5]),
        .s_axis_b_tdata(out_acc_6),
        .m_axis_result_tvalid(tvalid_res_add_fb[5]),
        .m_axis_result_tdata(res_add_fb_6)
    );
    
    floating_point_add_non_blocking m7_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[6]),
        .s_axis_a_tdata(res_mult_fb_7),
        .s_axis_b_tvalid(tvalid_out_acc[6]),
        .s_axis_b_tdata(out_acc_7),
        .m_axis_result_tvalid(tvalid_res_add_fb[6]),
        .m_axis_result_tdata(res_add_fb_7)
    );
    
    floating_point_add_non_blocking m8_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[7]),
        .s_axis_a_tdata(res_mult_fb_8),
        .s_axis_b_tvalid(tvalid_out_acc[7]),
        .s_axis_b_tdata(out_acc_8),
        .m_axis_result_tvalid(tvalid_res_add_fb[7]),
        .m_axis_result_tdata(res_add_fb_8)
    );
    
    floating_point_add_non_blocking m9_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[8]),
        .s_axis_a_tdata(res_mult_fb_9),
        .s_axis_b_tvalid(tvalid_out_acc[8]),
        .s_axis_b_tdata(out_acc_9),
        .m_axis_result_tvalid(tvalid_res_add_fb[8]),
        .m_axis_result_tdata(res_add_fb_9)
    );
    
    floating_point_add_non_blocking m10_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[9]),
        .s_axis_a_tdata(res_mult_fb_10),
        .s_axis_b_tvalid(tvalid_out_acc[9]),
        .s_axis_b_tdata(out_acc_10),
        .m_axis_result_tvalid(tvalid_res_add_fb[9]),
        .m_axis_result_tdata(res_add_fb_10)
    );
    
    floating_point_add_non_blocking m11_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[10]),
        .s_axis_a_tdata(res_mult_fb_11),
        .s_axis_b_tvalid(tvalid_out_acc[10]),
        .s_axis_b_tdata(out_acc_11),
        .m_axis_result_tvalid(tvalid_res_add_fb[10]),
        .m_axis_result_tdata(res_add_fb_11)
    );
    
    floating_point_add_non_blocking m12_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[11]),
        .s_axis_a_tdata(res_mult_fb_12),
        .s_axis_b_tvalid(tvalid_out_acc[11]),
        .s_axis_b_tdata(out_acc_12),
        .m_axis_result_tvalid(tvalid_res_add_fb[11]),
        .m_axis_result_tdata(res_add_fb_12)
    );
    
    floating_point_add_non_blocking m13_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[12]),
        .s_axis_a_tdata(res_mult_fb_13),
        .s_axis_b_tvalid(tvalid_out_acc[12]),
        .s_axis_b_tdata(out_acc_13),
        .m_axis_result_tvalid(tvalid_res_add_fb[12]),
        .m_axis_result_tdata(res_add_fb_13)
    );
    
    floating_point_add_non_blocking m14_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[13]),
        .s_axis_a_tdata(res_mult_fb_14),
        .s_axis_b_tvalid(tvalid_out_acc[13]),
        .s_axis_b_tdata(out_acc_14),
        .m_axis_result_tvalid(tvalid_res_add_fb[13]),
        .m_axis_result_tdata(res_add_fb_14)
    );
    
    floating_point_add_non_blocking m15_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[14]),
        .s_axis_a_tdata(res_mult_fb_15),
        .s_axis_b_tvalid(tvalid_out_acc[14]),
        .s_axis_b_tdata(out_acc_15),
        .m_axis_result_tvalid(tvalid_res_add_fb[14]),
        .m_axis_result_tdata(res_add_fb_15)
    );
    
    floating_point_add_non_blocking m16_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[15]),
        .s_axis_a_tdata(res_mult_fb_16),
        .s_axis_b_tvalid(tvalid_out_acc[15]),
        .s_axis_b_tdata(out_acc_16),
        .m_axis_result_tvalid(tvalid_res_add_fb[15]),
        .m_axis_result_tdata(res_add_fb_16)
    );
    
    floating_point_add_non_blocking m17_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[16]),
        .s_axis_a_tdata(res_mult_fb_17),
        .s_axis_b_tvalid(tvalid_out_acc[16]),
        .s_axis_b_tdata(out_acc_17),
        .m_axis_result_tvalid(tvalid_res_add_fb[16]),
        .m_axis_result_tdata(res_add_fb_17)
    );
    
    floating_point_add_non_blocking m18_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[17]),
        .s_axis_a_tdata(res_mult_fb_18),
        .s_axis_b_tvalid(tvalid_out_acc[17]),
        .s_axis_b_tdata(out_acc_18),
        .m_axis_result_tvalid(tvalid_res_add_fb[17]),
        .m_axis_result_tdata(res_add_fb_18)
    );
    
    floating_point_add_non_blocking m19_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[18]),
        .s_axis_a_tdata(res_mult_fb_19),
        .s_axis_b_tvalid(tvalid_out_acc[18]),
        .s_axis_b_tdata(out_acc_19),
        .m_axis_result_tvalid(tvalid_res_add_fb[18]),
        .m_axis_result_tdata(res_add_fb_19)
    );
    
    floating_point_add_non_blocking m20_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[19]),
        .s_axis_a_tdata(res_mult_fb_20),
        .s_axis_b_tvalid(tvalid_out_acc[19]),
        .s_axis_b_tdata(out_acc_20),
        .m_axis_result_tvalid(tvalid_res_add_fb[19]),
        .m_axis_result_tdata(res_add_fb_20)
    );
    
    floating_point_add_non_blocking m21_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[20]),
        .s_axis_a_tdata(res_mult_fb_21),
        .s_axis_b_tvalid(tvalid_out_acc[20]),
        .s_axis_b_tdata(out_acc_21),
        .m_axis_result_tvalid(tvalid_res_add_fb[20]),
        .m_axis_result_tdata(res_add_fb_21)
    );
    
    floating_point_add_non_blocking m22_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[21]),
        .s_axis_a_tdata(res_mult_fb_22),
        .s_axis_b_tvalid(tvalid_out_acc[21]),
        .s_axis_b_tdata(out_acc_22),
        .m_axis_result_tvalid(tvalid_res_add_fb[21]),
        .m_axis_result_tdata(res_add_fb_22)
    );
    
    floating_point_add_non_blocking m23_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[22]),
        .s_axis_a_tdata(res_mult_fb_23),
        .s_axis_b_tvalid(tvalid_out_acc[22]),
        .s_axis_b_tdata(out_acc_23),
        .m_axis_result_tvalid(tvalid_res_add_fb[22]),
        .m_axis_result_tdata(res_add_fb_23)
    );
    
    floating_point_add_non_blocking m24_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[23]),
        .s_axis_a_tdata(res_mult_fb_24),
        .s_axis_b_tvalid(tvalid_out_acc[23]),
        .s_axis_b_tdata(out_acc_24),
        .m_axis_result_tvalid(tvalid_res_add_fb[23]),
        .m_axis_result_tdata(res_add_fb_24)
    );
    
    floating_point_add_non_blocking m25_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[24]),
        .s_axis_a_tdata(res_mult_fb_25),
        .s_axis_b_tvalid(tvalid_out_acc[24]),
        .s_axis_b_tdata(out_acc_25),
        .m_axis_result_tvalid(tvalid_res_add_fb[24]),
        .m_axis_result_tdata(res_add_fb_25)
    );
    
    floating_point_add_non_blocking m26_add_fb (
        .s_axis_a_tvalid(tvalid_res_mult_fb[25]),
        .s_axis_a_tdata(res_mult_fb_26),
        .s_axis_b_tvalid(tvalid_out_acc[25]),
        .s_axis_b_tdata(out_acc_26),
        .m_axis_result_tvalid(tvalid_res_add_fb[25]),
        .m_axis_result_tdata(res_add_fb_26)
    );
    
    always@(posedge clk) begin
    
        powspectr_temp <= powspectr;
        tvalid_powspectr_temp <= tvalid_powspectr;
        
        if (tvalid_powspectr) begin
            tvalid_reg_fb <= 26'b11111111111111111111111111;
            reg_fb_1 <= filter_banks_1[ind];
            reg_fb_2 <= filter_banks_2[ind];
            reg_fb_3 <= filter_banks_3[ind];
            reg_fb_4 <= filter_banks_4[ind];
            reg_fb_5 <= filter_banks_5[ind];
            reg_fb_6 <= filter_banks_6[ind];
            reg_fb_7 <= filter_banks_7[ind];
            reg_fb_8 <= filter_banks_8[ind];
            reg_fb_9 <= filter_banks_9[ind];
            reg_fb_10 <= filter_banks_10[ind];
            reg_fb_11 <= filter_banks_11[ind];
            reg_fb_12 <= filter_banks_12[ind];
            reg_fb_13 <= filter_banks_13[ind];
            reg_fb_14 <= filter_banks_14[ind];
            reg_fb_15 <= filter_banks_15[ind];
            reg_fb_16 <= filter_banks_16[ind];
            reg_fb_17 <= filter_banks_17[ind];
            reg_fb_18 <= filter_banks_18[ind];
            reg_fb_19 <= filter_banks_19[ind];
            reg_fb_20 <= filter_banks_20[ind];
            reg_fb_21 <= filter_banks_21[ind];
            reg_fb_22 <= filter_banks_22[ind];
            reg_fb_23 <= filter_banks_23[ind];
            reg_fb_24 <= filter_banks_24[ind];
            reg_fb_25 <= filter_banks_25[ind];
            reg_fb_26 <= filter_banks_26[ind];
            
            out_acc_1 <= res_add_fb_1;
            out_acc_2 <= res_add_fb_2;
            out_acc_3 <= res_add_fb_3;
            out_acc_4 <= res_add_fb_4;
            out_acc_5 <= res_add_fb_5;
            out_acc_6 <= res_add_fb_6;
            out_acc_7 <= res_add_fb_7;
            out_acc_8 <= res_add_fb_8;
            out_acc_9 <= res_add_fb_9;
            out_acc_10 <= res_add_fb_10;
            out_acc_11 <= res_add_fb_11;
            out_acc_12 <= res_add_fb_12;
            out_acc_13 <= res_add_fb_13;
            out_acc_14 <= res_add_fb_14;
            out_acc_15 <= res_add_fb_15;
            out_acc_16 <= res_add_fb_16;
            out_acc_17 <= res_add_fb_17;
            out_acc_18 <= res_add_fb_18;
            out_acc_19 <= res_add_fb_19;
            out_acc_20 <= res_add_fb_20;
            out_acc_21 <= res_add_fb_21;
            out_acc_22 <= res_add_fb_22;
            out_acc_23 <= res_add_fb_23;
            out_acc_24 <= res_add_fb_24;
            out_acc_25 <= res_add_fb_25;
            out_acc_26 <= res_add_fb_26;
            
            ind <= ind + 1;
        end
        else begin
            tvalid_reg_fb <= 26'b00000000000000000000000000;
            reg_fb_1 <= 32'h00000000;
            reg_fb_2 <= 32'h00000000;
            reg_fb_3 <= 32'h00000000;
            reg_fb_4 <= 32'h00000000;
            reg_fb_5 <= 32'h00000000;
            reg_fb_6 <= 32'h00000000;
            reg_fb_7 <= 32'h00000000;
            reg_fb_8 <= 32'h00000000;
            reg_fb_9 <= 32'h00000000;
            reg_fb_10 <= 32'h00000000;
            reg_fb_11 <= 32'h00000000;
            reg_fb_12 <= 32'h00000000;
            reg_fb_13 <= 32'h00000000;
            reg_fb_14 <= 32'h00000000;
            reg_fb_15 <= 32'h00000000;
            reg_fb_16 <= 32'h00000000;
            reg_fb_17 <= 32'h00000000;
            reg_fb_18 <= 32'h00000000;
            reg_fb_19 <= 32'h00000000;
            reg_fb_20 <= 32'h00000000;
            reg_fb_21 <= 32'h00000000;
            reg_fb_22 <= 32'h00000000;
            reg_fb_23 <= 32'h00000000;
            reg_fb_24 <= 32'h00000000;
            reg_fb_25 <= 32'h00000000;
            reg_fb_26 <= 32'h00000000;
            
            out_acc_1 <= 32'h00000000;
            out_acc_2 <= 32'h00000000;
            out_acc_3 <= 32'h00000000;
            out_acc_4 <= 32'h00000000;
            out_acc_5 <= 32'h00000000;
            out_acc_6 <= 32'h00000000;
            out_acc_7 <= 32'h00000000;
            out_acc_8 <= 32'h00000000;
            out_acc_9 <= 32'h00000000;
            out_acc_10 <= 32'h00000000;
            out_acc_11 <= 32'h00000000;
            out_acc_12 <= 32'h00000000;
            out_acc_13 <= 32'h00000000;
            out_acc_14 <= 32'h00000000;
            out_acc_15 <= 32'h00000000;
            out_acc_16 <= 32'h00000000;
            out_acc_17 <= 32'h00000000;
            out_acc_18 <= 32'h00000000;
            out_acc_19 <= 32'h00000000;
            out_acc_20 <= 32'h00000000;
            out_acc_21 <= 32'h00000000;
            out_acc_22 <= 32'h00000000;
            out_acc_23 <= 32'h00000000;
            out_acc_24 <= 32'h00000000;
            out_acc_25 <= 32'h00000000;
            out_acc_26 <= 32'h00000000;
            
            ind = 0;
        end
        
        tvalid_out_acc <= tvalid_res_mult_fb;
        
        if (!tvalid_powspectr_temp) begin
            if (cnt_feat < 27) begin
                cnt_feat <= cnt_feat + 1;
                if (cnt_feat == 1) begin
                    feat_filterbanks <= fbank_1_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 2) begin
                    feat_filterbanks <= fbank_2_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 3) begin
                    feat_filterbanks <= fbank_3_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 4) begin
                    feat_filterbanks <= fbank_4_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 5) begin
                    feat_filterbanks <= fbank_5_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 6) begin
                    feat_filterbanks <= fbank_6_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 7) begin
                    feat_filterbanks <= fbank_7_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 8) begin
                    feat_filterbanks <= fbank_8_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 9) begin
                    feat_filterbanks <= fbank_9_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 10) begin
                    feat_filterbanks <= fbank_10_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 11) begin
                    feat_filterbanks <= fbank_11_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 12) begin
                    feat_filterbanks <= fbank_12_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 13) begin
                    feat_filterbanks <= fbank_13_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 14) begin
                    feat_filterbanks <= fbank_14_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 15) begin
                    feat_filterbanks <= fbank_15_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 16) begin
                    feat_filterbanks <= fbank_16_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 17) begin
                    feat_filterbanks <= fbank_17_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 18) begin
                    feat_filterbanks <= fbank_18_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 19) begin
                    feat_filterbanks <= fbank_19_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 20) begin
                    feat_filterbanks <= fbank_20_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 21) begin
                    feat_filterbanks <= fbank_21_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 22) begin
                    feat_filterbanks <= fbank_22_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 23) begin
                    feat_filterbanks <= fbank_23_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 24) begin
                    feat_filterbanks <= fbank_24_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 25) begin
                    feat_filterbanks <= fbank_25_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
                else if (cnt_feat == 26) begin
                    feat_filterbanks <= fbank_26_temp;
                    tvalid_feat_filterbanks <= 1'b1;
                end
            end
            else begin
                feat_filterbanks <= 32'h3f800000;
                tvalid_feat_filterbanks <= 1'b0;
            end
        end
        else begin
            cnt_feat <= 0;
        end
        
    end
    
    always@(negedge tvalid_powspectr) begin
    
        // ���������� �������� �������� �� 0
        fbank_1_temp <= out_acc_1;
        fbank_2_temp <= out_acc_2;
        fbank_3_temp <= out_acc_3;
        fbank_4_temp <= out_acc_4;
        fbank_5_temp <= out_acc_5;
        fbank_6_temp <= out_acc_6;
        fbank_7_temp <= out_acc_7;
        fbank_8_temp <= out_acc_8;
        fbank_9_temp <= out_acc_9;
        fbank_10_temp <= out_acc_10;
        fbank_11_temp <= out_acc_11;
        fbank_12_temp <= out_acc_12;
        fbank_13_temp <= out_acc_13;
        fbank_14_temp <= out_acc_14;
        fbank_15_temp <= out_acc_15;
        fbank_16_temp <= out_acc_16;
        fbank_17_temp <= out_acc_17;
        fbank_18_temp <= out_acc_18;
        fbank_19_temp <= out_acc_19;
        fbank_20_temp <= out_acc_20;
        fbank_21_temp <= out_acc_21;
        fbank_22_temp <= out_acc_22;
        fbank_23_temp <= out_acc_23;
        fbank_24_temp <= out_acc_24;
        fbank_25_temp <= out_acc_25;
        fbank_26_temp <= out_acc_26;
        
    end
   
endmodule
