`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pVSB1fdp0d8mtg3LHrLYCqADYNQv1kYsGBMv/+K08aLxh/NLENzMM7hXXYld+2Mgd7vecGpdaC3k
gwoJ87eJgg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TrvLQEi/uJPAZXHsPaV57yoJ9EtvRVNbWErIxN3rJpRzIiClrcH6SWry1U/juttM6Ef9Hp5zSiEl
xNpXxoS8wD1iGQC3wTWm6onL4lbs5dCr5r6SHKI+yRvk7PM0lNGSuxzJxiESo15OD+VI4TBDw4Zt
hcxOQOC9HXnv4RekyhM=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g55PFOQz5gBNNuoAKJA6LG+Go3evy8K7bR71fr18lbAHBy6BXY5cxyMVmR6iMXA9xjvLNX9ZwFxL
yW9jhdIKz+0phA20qrgB9zIyJLsPj7lBLFXWAKf8rmqv2GMRf7GqCtYK5Pqn6bxMwn+n8j50ca2O
X49Iq1oj34Zh+mics+4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JjYKvrh9MOLSA4mR//LjTlBGaa8xCFhn+/gMizL6ZibhVKAfMan42h7Ih/5YTGi++UTn0LHd9NL2
NaEQm2v4o2/CYXMF02K83EGT2I0yUSTUGc3tcxpNAxg390x/Pf1S4xXOwpqZAYLjhWse/4qzYHFe
iIQp1rnWICwKmFo+ZDG7yZ46pqq5zbSoc4y2p8g2Be/9TN+Y61xI7+D+EAu7QTdwsL8a3QMsB7Zo
r8bdBBswbfd/oqL9KLKL/Se74397O2HGv16SR7618OwhGC/PJGF62sCa/WzAZbXDjbk7bTLUCyoY
71dLV9qD6596pGntd7mPSMKPXsrBqm2dF4MJ1A==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SSijEQc3z4IgPRpOXyZNPGTBKNNDh8UIUp6Jc6nCd2BhqaRyKvYRVaSbO28FxPLannTOttVNc7kk
nl077g777DPyzXTsDcYVVSgCq66KzFzd9air6Rm4YQEnULnroQEEBvsGlrlRApzIY13fCR8Q8Fes
8flh0wIvt1IUA60/FMM3YwNPai5m3k19RaY/qsBdtTNLM+8XqaS0XCHWnyA2QHtb6iqRTQyHXNpO
tBGXOMyVMkyGUq2FAx9nYlTvIbXYYvrUtsQaGxetWks9vlDulbTRAnCFb7GU0+h3l3y+hF4Wzkn2
o2p95CyRx1FQ/Rn0oxBn++Rtk6p7bYPQS42cSQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L337KT5q53NKw85qdeX1tBHCmb9rh0WndWsKzAyylJ7jXE+LkDsZ1dyUX2YUpfCn9BKLEH2MzATq
tqzbaiVWOu/xeMRiU5/wkXL4qEX/dKjPRSJlNBWwDa9lFGbdFy89cWFoNvS+Teu59m5yiiDnIsEO
MXDu8nBP5UasM+BEuesC1UlPIu7vinDhIbxmSZZQfdQoxRJrJhS5MUcMYRs6Q8mNJvPXbo1WhUGq
lCkeJ1Mwf+GUzVwd087Tb7Hf3TsU6tjTfAyqJFoofzOBAnyD237xgkHu2B+/4AT6bby5CbEp5ISZ
1Crn+G5ARbRRqoqaFdx72snFnkZFJIffkdR3DQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 119648)
`protect data_block
3U+9z3xqvHNIcHJ4qx56r/rIXlWVfpX5x/9mz2LdIe45MyKdNSwZ5H9ekgVHHKw54QTFO+QMIKtL
nrdJO5883lCy5qoQpDBO1IkgJtf2q7igNxz2tgddfHwQXzR54FYcFI2jXT10ikQ5JBQiImf0Xbbw
Z+qguy2aj91LStucA8YJSEUtOOKhtvvec05RcCsZ10RTmBlO1+E0VsAs0VCRkAAYTTD+PNy/CG9e
QNWSMzGor9fnew0IG58vLn0/O9xPbxaqMmjVDuTnKaWU5mDzPwV34yQ48hr1DMDS9Do4oFDYjkRw
f/Aay7BSb6+OOh2tWkvbdilPf0xk4tUey3Nk76kLLgVx31lUzi/jBki9Hva2DDIwXEWmZvHP4AaC
5pzeXUVTV/mP8k19g/5sP31tUBIIb1ZcGem+KDGS85goCFHNODEEp70WfIJpo3eZvNxJt++XBjGu
ZheVWcnXoQE7wc+84Ti7y1IVFgwqS9XUpHtQbqmuPsQLHtAe+9XHn7upEGdlQTkZ2V5UEJtAAeqM
ZCuOO0aaLmTqi/+Kreq46T+rdXDj30lmfZ+5Bdx2QsizPIwUAHsxY9Z1O5cM8eyMkbI9F+eqChqn
TbiWskJRn60JCZ93CVH0Ps+CJ5XPrNBlDlJ7ycoNEqXZtvbv66Ue12Rd2J0ohMLISMUe22pOFBfr
K+lRcA+ZLPiE9qBrGbb3qh502hrmuAOt5YQZdCrgrxCNtj8vqmxla57pGLKjzzff6gryM+JAqlkW
Y4Ew/D44GFAHxmyygVV454v0K8NcB6NV1cEssXMfL02rCr21EljwTrXw07OTEotRwJykYO8G2LzB
xJGYW3E431M19JYe2rLPkq4o4e9lpCNHWx/MnC2zQWqztYmykGazLNeikoMI9EPXyEdaUqMN4tYf
ipyGV3c97kxBUBTWUnbpR6/xXD4MSm0jVdFl/TIgZn6Q/AtuRJApVfs1ijx8fM6dDm6F6xSN7ez2
vwB5IKpxqyUsm0GWD4jtkx/2SUgvHZJ0MvvP2qLfTVlJhCYi5SPVfhtHg5vfTmZjVMaocRbSTC99
4FUgHnVqYDI0AtVvepC09UtaPMb6OM4uh3M/8ayDkFaHnn/bUJ9HlSRBE99fgec/22S8v05xI44u
K9uw3wVXdapJPuXjzF912vpWB1dhkK9+GfLi7hq5LH26AleyqmUxq/niUs+oLwlHfOKn0thQNHfo
uC7lnPjzu70gKBlkqgeVzW3AefrqsksYABs6v9OssHHkcJ62pdbJWW3vg60MgshFWZyog5+RpOPx
eFBmYin4kJNJ/f4F3CdvpiIrCB4sTLLBNND4CgauokZ3PwIMNxyQ3qAPswq0OG/XT8IpYxBE0w2c
siSDHcppjFcGnObheARPnzDCMEwwrKGhdTf8UxWjqliYC/RMAgWF4sxwAYt46cVl56gqL9FFa1TX
I1H1affwWbbZqtZ7lj88noyW9dj17PJzRGQfhENMbUicEakVoOmFMwuAcD/GUSYc9qsyPriLInYq
uP3e9YVkYuNgQrzXZEmcpObf7fKQsGKkp3/fcDX6ZIBwV/gzKq5kdoHzoZkqjD7FuzzdVVoQfWFo
lomIJpCGxU7N8aR9tCNZaQxR5FiYWF3Nva4IL9ykgONWp4Y/VcVslM541unPdVl1/Gn+9dBGv8za
8v2v/oFkvOz2ZH8H6/cadJjwfGgEvN1YzdC21Of7BG+fBZe+7KIAN6oA4pVdkxhMjN2/nXKum+H4
6KcGMlvTfQaf+zh+Sz8cGIP0DgtHmQ5+uFoZ0sN9NI9PN49Iad47g6neyllTjMay1FJHG88aGO9S
Ef9rjtLX8LeokKLCm+ZYdPDnz01hErbgp3GVS0NnJPoCqFLi6p8SvhQgYJ1XPzD0dMeTyUlx8XX8
+2o668+qIM1aV3saoEMmLRz7QOAqLivYzvNBww2mmw0qvdeiJsF1CTcV6eenIuXifveUZKfA+SgR
nEq8YtG/g55oUbAQu+3IdRCNWigYW4OsfzQoHiaD3AZxiWbTQQcbhuUKVshKeILfyR8zaQuJK00X
lXkjDHTEev84OxusPfX3gy3Foeapi/Mh2iO1LMDJGMy1S9pl/uNUV8GXf1O/MDlRmPGEE4mIEgZ7
PYJl5LldhiePTM0E2mHq8zm9W0F+0cFOKVdFE5UgVrUmnVvGwRLEvNiWUu17eTCUUFrFEOfZZjDc
j3pI86UZyB6lmcfujW4jt7YZpyfgLgm49i0BsOmygO0c55xusAq/8f6FApIanH0dAFoI9FScwC1e
4jvv1BXOwfFGS8hyg62bYoc4zhq3S52fcLIa/nBgWcE6Hixyk00kG1hlH718XjPRhGt3vSgPyU5D
pdIi/G7zV217V6slhXERxE9ml2Ch/DO9iLlNVMVct6GOCUfei8wwQ459eoaqU2T7a5mnogjiUd0P
EfMcqD4UZQZmOHNfkCouOSstdVqCEzBHCchd9EI+6fW4Rfc3xcuxS5Ewq35CoHdQ2GuDKv9X+Ba3
Mwt4ZI1PaxJIpfPKNwjtQyv+SviVc3lEMsPy8lvZL0r/8jdcmpkUxIyXTetA4f48C24eBPDMYObK
dROmvAS6Ip9wx/fk+trzGTFzpc6tOUm+WWkAERdrlA8JI7uhsKeJ5DkHhWXYgOsVe/eUHuXS62UZ
UuLGEINocPw7qcnqEMGHVKOsN0BsO4OTmOF2D8OdFWBg4oM4UPIOvpxPlEWxhZOf6HnZ3RE9CNBC
DXg0+gtft/iIdMjpZrSYgGHm850pXDrOpiMM0YWfh/3SkSFuxJuPgamVUA5fof+Qvr20P5SlA1yu
Qf5qf4BlUF8y7U9/4XkVlTFNLIciC57PdgtZUu9DwATse30zIYueYvZfEofZHuWCNzf/ez6DVc2V
F2ZUfR/3fWprz5cmfrCnLxA0xsyqWHSHQfazTc+thawG8ff9vIU+XV3HY0qTvGPYm2/MlheAJEvt
B8NA8buo/ydFwlooaWeUe20p6PtyRJV6vNzbOiWAhYw1uOeEmzw31iqJm8rSOWS5iQBCw1YrPb+S
AVX9HmWLFW4FVSUdd4UiuF0KBuS0VhsFeqU+Lz9B3HhXZeRvBYcYm9kDTq8sfdrD3vtlre6b3SNo
FXUA1kLmWOhFH3FQDZ9oRYN7YZ7rpNJPBXw9PIthHDJujI5iLbKZhutyJUG6N/2/XLSx/qfXoWk9
OfudwrBa3Fs0JjsxB/UxlNAicEmsrJZ9J4++CPl9ETVgHLh108ojE+/DWjtvdZMcnz9SJ8WxKFNs
L6L8US+jX4rMd2l+psqG3PJuI7LS90qdn5EpPD0RXWB/lyVQgyGAA5cQYe29rfPqcXBD3iWDYxcD
9/ip3k7ZJa8mDt49n580W75MAffhLLSPsNGerDbJ86KNZiz3w9a2FcKc79r7qA4jLHUQY4+OOELZ
/cmAKoMuR4SWNfvjT2V/bii/W9Aa797NzQg18uqKRH4O3M8VtLtCGxUfjrpOiDe4F19uz21tomjP
z0xlwatjVBiysQ2DASJZeCFCzI93wCVYiExHBkM2PSn1D3hEmQMlVP4MDgEf3t4diEsOjAsbKuDS
RdoxD7bN5yU1ntwEE2wx2eLCpc5e5E1IMZFYQ0wCyNuMVMGWpwzhpKy06iG3XDxLwG7diB3PoTql
BC9nEo1anp9FfumYXwUb8/b2JzUCkdalLhUXMgv8xawCM1BDf79DxOo9r0llsvpaPXciJ3KbGyPb
uTW5dF/MkZNeT1eLRi3mv6qKUGaa28uSxFZ0GCpsiw7FYY9LAhNppq9n3Abnj4LQcjbKszmcyeIa
DL+eHR0qZiz5VOGPQdqaSEMCDGUaK6Ir122+OFAgIVC5mLh1UInwyMBXPcSPV40pht+2aV6aqxhW
qkk5Bi3QKipLe8BO/qoSxi5o3eMlQZWibqlQLX0Bv30a9Xl4jEw5f6hqfQoimqvdx1uEVzrzuSjF
qThn82tmaAKvBs9dMKkqOMCvX9pHGIy8759kpo0mTJKb0Vk532E8J32mVVs1yBQbNXYuztQJ9qjn
hr3kH16fi4ZABeD/FNiDkOvZ1rDVUgYMCu5ECMLtv1iei6DFOsKyDm/vOHNqFP1mps5szvC3eYBZ
CTUzIbdLTwYrEf8B1Vg9VTEF1hAEf7RvX5OCRl1p9Tku3b4Pl6W9E/O5pQ6QsSXeIJK6jOP92tbr
xvmJi700GFQMum63p+inGTFCYa1zTO/Zyzcnn3wPE/Kyn64T/86Y98DNNTc1/7H1V0Okj3roTuXF
RSqNwUlH8CkuOa770eAoKonVdn11tFaAVfJ4e62hPVUlpEoZyfhPvAgGX8KaQjX/nwBTEj0Ptr45
ukaIWnHkiU+YCUK5ZfFLglOSM4lXyLdejBBZBqQcJl356d+U7IFMzmS5MW83WT/2taoy7QaPLeUm
Q5oWDCjrznV27CLKFEHbTEDNHytlJDTzHGJpMNamGl53aHTGEF4D1BLVODUUD0ddvIJt//hsqyYp
QghGWu8kKsJzM9PxJ8EvFCjPSlQHNeJ6hfmK5D3jn32gxAw3qblq3PZ6zgnssZWvmuyTSjPLT2GP
2I8fu4xEYlKKkGW9dIHYYnK++Bvh8wseEJYxFB93ZPYnAFS3RtHGJAdQn1W9fAeH000PELqgib9+
2EgVZhG/iyKCq10/Lbex7jJ2zVvmtQVoijWOu2F36aEy5NOdm9/SUe8MqTyXfhOswSpsfvQmmgwY
pe4qIsmZG2FD8LOs4+i3jKU1QZuf8baKvQ4EMvMZYfVyB0M/fe8ngd8ztEwbERJbuYnOejjGxiDo
br3Pimo+2NVrh9aGsmTS0XLnNFsxL7vVn9fDHJGMehNn+pke9G0+QWQuNZi+dVGv95q0UoLHoXAO
uvVgUvPJvYhWNfeV4+gNsxqdlNUisW3ETFJP522fSxI6Drwigrijq8g4TVNSaYns8e0ed25GMvnW
Fz7u6KCI8up4rxV0YC1Xw0snyZ3NCONAtZyfgzYWI59yf9DpNLaAzI4U5kMaVzSRZ9SpSM+bebyq
HpmjcBnhBQEVR7Szhs9OTcZbIMMatqW1Q6dOiTHTZNQPqyEZeJ9ez+7Ov9ndGpG4gj0qBZUV6SKY
nELVZzEHtD9suKRamGKMHfpGixebGYcMGqAflzhtk/JHHrz4GRej141jdvV9gtnfNptpdzcn2mLE
aBL9rRTmqVg+c7Y2PRIfJsrckj5gaG/sAxMmNVVkjEDQrJTJsyC0A2ERw1ByIsg69GiJ72+EGIAa
TD23/qzOmfAh6BIzWYYhgOYbuft2Dis1UZPj39cJpYbf+W7M/Q2JGhYu3hFMyExAIdMeNPldV8gi
h6eKUsbE0COHWmu+mnJFsFoMUXtVSIm2se291jYwcaBLv8z1gg9IHzO+5KhImF8J6nKADXZjYQLl
r3/O+Ra/DJ8E9fltnwqcPiQrogZd+pBl0jm1UpAV0XNeBFzVA6EjQV50mRQblpO2cucTK/hd4kv6
NQcfbpmn9tHOVZ6ShZix4AKAVpZp/cgv0jTOkulfomS8PouuY2PFJ9mwGMtSHfczUOFJVKjohby0
KwbDtc8Pj75o9QShmxX4DijfQFMBrny66QyDaGMiYnLnICwR50NipVX+8wgXlsPhdp1tqUUHPflY
zLTeB7hJDAa+LvNXAaBeWtQImDrbXQc0Tq8du0eaLAxd05VYz1Sg2+JbO9YYXe2Lx/6y0NoUT8i8
QylVGFP6tjvhS5nvK1dp85gatJ+6UiOyaXXWCVkdY9R6kkgIun3sX5YjGhoduTjFh9LWhFXfk6/5
OxEgGNgwikHhpPDMV7lwiFU0SbsOS1XbrwaT3J+DsW//grQ3aa4nCcbzSZfrRrpo1Jru3IAl0gFw
xw9lbbEd7aUjClVCkfTWXqFyL3ApSANZ79HqKFtAd+gWvnGCpRomnIUnnZsTdfplEbiSHYenePtw
vTILRegzkZoMqj6b1nVGzwiaS/ikpdb1RBTvt/XDRr7Qt67XDIN8VhyWG5EvpL0vubhc4MeCcKKh
/VhsFqdKvZyVacv46I2JicUMNwjvYHsqwIhE6z0i3rcgxAe3fN0U9p8MOORcYQfCdR66CbMhg5N7
iUwYrT6mZ7U7PofSSLj/afbowyaGV7KuH29qJrApe1prV1FF3qPs2oMe990IxvYnDYIwFlNWwa/y
PhRPVHEAY41DPc2Aazuu74vz66r27oQv0VlfpwMhDKdDGicbFObLQ83Bxf0oecpCHekh4vRjpI3Y
RpsJEvljB+3tf4c5jtf+nsuAFXIuWU7HaWmpCaifdW8Jq7f7neLwzvTzHFXZw7WPWQi12R+Ylvif
mMLT4Nr0jyQ4QGTbiPgyJCPOFcQt/pMT3GUcia0maT45TkKo2Z1QmC45z+T3ESPq6kwqp7IiRXvh
RDMjZhJnPRgKGBvQKWIljqQUo0tj2mxr/pn7ocZ4tZIvX2rTl1RDaatQI0mLfUPWUUqB5tF1DYK9
k9i6sh33wFlDKHSo30T2LRm8ra597XRjepCQeOgpul9qOwdf3trDzDyFpfsUf41fBYuNcX1aysTL
UwEPa4DTn25j/XXgcviukb86GCIPItny3bbatlnTrp2PVXqmUEjfcISPo+8zY1BWaJdK4u5ihPeK
+Pp5t2GoNkjwt/ITYVu4pbThCAvuxVSFQnqmBOggXC42qdUGEHPuV5yZRdodHmBzdPa3I1Xpj7ts
90Mi1FbyJaxS1xK5yxK9/bEU6t/13MxWoIEwNUWATeac+oh983EjfEEdDGK5zBetcx9rAakgjha9
M6WVGxsgZcckwBsB2/cHOdKFCnmmiYK89jqXIXPz/HNnFdMjhDj8WfkDoMCdSTYq+go4izMHq//s
/J1inntwY1fgBvoG9r4ehxM4Mamb2FmEst2CCIrZ/jlTufIemyuCjf/Kd5TMEJF8uk5QBxWS0Ohl
EMcIKS8w5Hsoxzb/FqSkiHrtjSEZMbelD+lMcLKe8CxtncM/1j70BgVI1kXIeaQYxgXuZXfAdJDo
3k88yABEXAwasb2PV+2i+pGKMymtNajxeUMUnDoGsKA3/R1jn8T4G43UNuHd9IOTVt3UThjOFYGz
TpcPLlLsufkffI1l0f7SuG1NaUQiFu3zXPtZi6IVgy7poPiJSEuj9vMbdo1sWs1E9tLMLH5UIE2s
gS4gMQ00TwHREboRGqH2MhYJP4YY51StCtrm+cqXnu6QaE4888g0CtwwIjI6quYPyY8hVrZZy/Sz
dXk+q0XQbvK/8JjUzb2TT5sWFwCnb0/+YYq0iZPmirNciEkNHseBciED6lBSS5DK8s3rA/wo/Wp3
InYz/Ws9hWvo4ZfZlUuQn08TdoDguqZGyWxB6sho/lhnWeFFMw2HRKhdAlyui/+v1Apf+RnFTSUz
Xp9MUzmeQquyW6T5zknmt7pfoGFuTXxOP32Z5ijbNgDevRRBXItR1Nblc+CEIHX6i0+mK8Gznd6i
Rv03c68TDsQam0VdfJ1PhlOriURESVp/W4O4/BosCcyYMAjOvx6IuJpWte90fbAG7LAK4uoXdhhq
tqZNTdc501eHL/7at0UvXgl3zbGsOugUw3zqk3kiWPrSy0/xNekWZuVxmscovjsjadyJwzOO7B79
Q1GKyCDE8dvCIZ5VxABkdV8kjWcfaTYI+o6umUVfo69sA4aUv2phQWxH9BcmnFhOA3hS/t2MapBd
nVJBgT5aTMiizNKNivuZWgLM6SN5QJePBJkB8jMXlyza+KPu1UYDf6usQju2V2+5jEJ0+xq/CKdB
ncXFMk+fxY1NzkCtbF+D4jmhrRQjduSxYd49BXqlCns7AZszaM3PL7Et4TcE2JHuJZQXP/6CzvP8
EBrXdxH7bBQtJdBJ79jKuXS9UZ7UJd5b5hlKXDam4SwKB+VGnfwDFPreKxrEQw1Ws5Ah1RYvpX4c
9SmLmaDSo59g69QvS17DDO1hfWkQ5GeEaZwCfOyIyzBXbvFxyaTXrXtPVTj4CGT96aL8rrfu0Uip
SHoSTfGeifCAYzrte1Xkr2n93Fidj1Z6cX7OYUAEgwF+qVOxTr/rKeIxbz4fe0fOp7JxcwsIMR03
c4nz0JOWYCdXifvQr1lPil3UKfKlI1FEbVvr9R3XOIo72VpI0UvpZBsSZnmzFrY9QEYzIWK/Iclr
rDnux1nuKPIJB6oLnokvshK5xDjpNTYTjwGFQr9oRN1w/cVEqf25xu9TqeyZdvUceA60j0saGzaY
WiCBEGcS1f8omsh6MzgSNKCKFZV3l273mPhNXY1v0GRXD8Gtt+Usq6yUrJKYQdT69Lk3ifP/kr/P
IyLZojYtJE9i0i5B0NGjEdx/wAzUde0i9W6ehk5xRgOTIElLcppSxA7pOrOCJrw7KKgAn1jzAXZh
5Lt6A24JSDbg46Lt0Cl0MJX/JNXPV5hKa2TaZzEDxZbH/Xy1xWXAuck6T9++g1gieIHsBVKIWUso
ItWlXqUrmJs1hGtN9vHW865lWfixnab02RnHDvM435H93egctpX+ZIq20kuOZwx4DM0BgJ8YEmVf
7d0i4qyCkMXnn7JLUdefU5GFWwtEuLDa64knrrQ6oN9WAyP/aGeVhYW4nOXbokbXNkHt+3F1vxU8
cO0kyMLo+l3P6Rjs9mYAYztPfGZSpLEUGjCH9YF3LC32ErBi3GIZCSOq1c9AidtilGtFOK28aYnk
XINzam+cW8fY2u9HFFBoRxWxtyE+2whxk2sLGD2yOy6Mojfh1Sy8fi237Dlo4m28yY3l3aEfxCLz
iWkBacHD8iz16wowK76g3hnXkBleIYcsaLbLO0Mp3/jPeOG+YJcfz1yEM/trXcv/S4Kn5ibDe4CE
3eeZ4UM/qJXmLntKhvlCRgWrdZ7AzUUGw6uj2KwHTxVyj+rru9BhyQcWsbcfTsxj9Rx26+a6dthW
nja6oWY0UF+PZYMtyX3qGYaNBe/tDVpXuywQgpx9LK4XTR15DoANBjNmkxTB19ZRIfCj2NrgIoq2
HWepwsmxz4fPazI8tHGCwFqu6EiKfRUZjiIzJPRakPp80TmNYmQ9VWFLBchPq4cwgTyxu6HeXRpm
GUjmZyrA1IEW1Af7tMNv8rJDXztl/XBUoT3q7oXVjB1SkwnkGMPAakiplxcpcoGDiE16vZ69EV1z
1Y8RYBNWeKgFDqXNuHyWz2aExzSFjp3HoGJO7Xdr0vQY7R+g5vwkFBULCGFJxqEcZueciIS5fxbM
q9H7G2ym4o3fJTTTAlY6+6KE6NqR5RI0fO8smbtsp55eWCPW5jeovPc65Sa54yGxWb8vYzZW4SHY
aEb8FIJFEeBw2GzbRlYBbtQaNsAbxUYR9HuBKS8+bx6UGwqBfXp0jsUddONyHv4zeX30rOIqIQvG
m7PdcSsCeKGX6gp6BvBV3GpjofPJv1mxah7ZiFzp8UI262g9WLe61gCQq2Ch3lpYjyZsZwt+BDuE
sy5H8fuiUFPuDYQxe2BeUQqzBNSaNYziMOYCpS0OWvSA27sdcjozsljji99sct28HG/TmCYikY3q
BiTGaYqeq0/NjK8wJ5oVGIgnH/WHYvieER8135e1yBSR+B6AU/k5Je60ymr6pnyIIlBa4e62WGLI
bfnbZY2qcRuQkGrraPQnYzk97NibCdG0JI7lebKLwVK9xAEYGBWju8WZtj3Hqmi6NAQ4nzL7WT14
9S3AHKmE655Ncl7ncF85qwPOY8tCv5Ko+EIaNoujd0wDKcxcMdqkBTfdftEUYHiZ6SzlXoQDhScV
rKBglA5GuBtAeD+aEhin8roXOoqEpm0s/azXdT1/FU8NmVsuInjU3FSHpAN64DKmVfAG7Ig4zgNs
29WPQMAS4xlAT/X7jFsbcqBwLTke2XYTyp6e5XHAMHWUWW/9OrTuwz7FfClTVcS0mduunyiBwgOS
nbZ+nextuMJsgAcx5JZTkf7a0hp2ZeXGpvJmrmIiUtLXw0xYKq7LI2dhznu9GORCQop+ZC1d6Geb
0kPCrGPpYdpQUPrtzrgCiUgTIUFeoK5LvK1xavIkzrCupUCvbwrfn/7/Z9kmTBbwTFTByOebnqQQ
3iG6Llr15EwNg6+NJGYQIwXEHJ+DjCCoUZ+yXLWBQA1TocOzAMktimIgJLx+vC9V4DtDHdM58xL0
n3j4I5mjNgj/1kSsmJpSU53mxYV7PgXtXi9dfUh0M6OjI63EI1Tupf1aWnuGzBt+J/QOyYro/GtU
OPO61Zv6jMVlmLmh/4aNUjdKuBdtBomPXGr+JWrqmgolhihEZ+Xu+SSHsVDJoiBGpAIwkQOn4GIY
qBv6atsGCcqcPqHIQc1rZD+WmRze5u2CpR6WRMu+ISH9qD37sR5dlNXJJ4DX7+/oReJA72cqMmKj
WNO98yfh8rkFvCrSSuXq+4RWNZIprUFjTCBHJfcHJy1fvmPavMK1HjvW4M3BHlMMjKsfMg8sV0dn
4nlXPYst4b1WSxfcrGoQk9oTZA8Io60AZkHnGDRtpwNVpBMOuBHEUipgVb9+Jk2qzPXgiLuCxZpg
HMR5z5n9wDkOSNxlWecf/j4Fehjhiz8LmA5ubNT06W+s9PNlNJRvGBdBgBxkieAFRyaqevZB/jlo
MfC1A5IDTogCcpt0DWNX6bt+YQMB0pDn1uK7nPg5AUntOf5hIj5q0+YeF4edrJVAvYTS8T4uFiPY
BBgBFHghhAn5ReGMl9UetTYYMfclAIQVUy9jZRbzkrpvy+6wZlcGkhnIh3t6QiO4dspR8OUlokLA
fpvD5aARsGxPwTfjXXDqmp7lnfcUJFPEtisyRAzUNXZ76e5cQbNU+Bbtz6sjnZqwmcFL054funpC
OHB/SRIqOTOp9ndgfyOt5NxE57lTxyqCHfIAaXG5XfnYdRWpgQ9Ou5IQXrCFkukz3vpwxA1QkYME
GOwf3Md1LyquN1VPvrLYx8bDPv6gYPVQss9jjI7CMZjhds4BSjNk5uHiuEgLCowqcK25G1+nJ7Wm
n150Me6Adpgx3Ir4V30bTBYG8T+kDW6LS02/fumjjU8CRbg3BYVqUXEdYvi5D3A7OOlKG98Y4z6K
wvTA+6ZgqWk1MAOnLd8X2owJjC/mbFqzQq0Aq857eD2x7Oaaiy1ta2hJdsfCH2udTBq/NytegPiW
MxIWEPqJfWsZqeYIrnjK8dRx+sM2MFS5vs+Gc1qgcc9WWeUHfzMILYlq80+Ru8hYJ4SltsvXews+
IHwNEIPDuMvUNgEwtXzanSAI/Ibsh08Iz3Lmsq/QrZUNb+bYTaFtEdyu/cOjA41GcQPgEEhqcoPa
6hyKTAHDnplxwaslPyIML89ioTL2iDW3SNSRsIrrhWWgLjHbaDfh2NrWFI1LpWHLgH/Y3yiRoY/t
L24EqbhG2IHNxiylArHvXD/fAb/hu8sUZxR1N9g+fm+JgBgmPira6m3DGCDHLsbhWpBP+g+DvLIe
9TibmqG/L2c420WrTtd/2FbHs6Zkpl0Oo05WH0uY3ZBvxCSO0IHYULpNk0Z+EsrTkGqMCOGjDMW/
km2F+6F1QIsqrF6yLDuYn02bdLzklAcVvH9h5WdeUbCNIDA9YtiMP7PiGqf1t6laE2VMseOnxJk9
Ez4ifehPEITSSf+Mj/h65teoRstBvbhoa8LHNZlvBGU6XDtdnqALcpfrqmPGUv/vaZy6T5hnBS0j
J0d5tXr2P5byWuyO21wEtwK1/N4QGDyRd/Dm9Omjvd1aQrGUVFK9EbKM+s+LGokbvJmNafKusNR5
k5XCt7A6sG3IFh+Gk9UQGO1Q7fzkH2pkU1LM1y0Rvips7DmihFlZj55ycUdgRzEzb/zdEoabPSa3
GE+wT4BHswntneHY6NOl1etA1fskOIpgo5nh274a4EYVpRLns3N880ef7xKHcPu09iDIsOER7j4u
JG/qzwPuoL2WeSg3XSR6cNQA57CJwtWxcv961aeG1xKr/XlweNcrgHEqG2BLBnDJ0bdU913VXyL/
kdtZjctlQQ3BTqB9oz0b+tBsb5TxArLMXi1A/ors2GBVE1ds/h3E7MgKggE2Ph/KDdXCh+L3x7S9
V4a8rrtlYOsOPcHkKy2XvBx8tKci0sL/Pop9F1A00S5IOPb67JwQSO4ZXchcQN1a/VGxD9587Uky
59A88OhEH9CMumlpw28XQFjVyIQ3B2prpctx5x6El7IL3RYBAtuNQDuhuXJEbmMHz3W+2SGKnqV3
l5B1kAi6L1qjR6KPK937gepDvkTPB4z4OspIXf2tUajWRyfCm+Upe9YAgmtOA2x3vsrcWttQUmYI
qJ1L6fSm2xPNRbMLxJJki9pIAicvUUB2wIUX1keQJsLxflLQ/XICc+T0+SMBHtukQTkEs7CIPYnI
uSQ4k0tvWwqOaALftN/14+nidkffiCUuErEsvDNndAaC+kl+JASkiJx9pFOWLmiQjci4zVc/B08T
YGHenvotcuiIehNqNP/JO5d/nG6fDdTAetkFBQ/cbyvY8XkT6PMpxvihda8JveBM3AjzHjGaK6UI
16vR9X4w41mnziHCdm1l3KbMafuhcYP/LbDPcbMAhqo3bToe4iLOyADIRa5A5FoOu36qX8vllJcN
EUp3mZxrqe7HQakN3+tWOHJzKbT3y9y78hukDlINvcHlEXTFCizDTCaRcQhcqxhx2URX0bvgakvk
uTuE84arSP/2vhFhAkOSjnpt7NeeGRK4kcZhW6l3/UJR0EGTbJSRrUeVT0MUBxpoYNJ3SgIt5bmT
j0YszXcL80wI7ppu/ZQ5kg4sbQCQ9A2TMa+8M9dofZdd1460Jer9E/fxCm3+ljX+k33pJkDEyo99
7zZuWLHQYE4vBXtpOi8c3lJMpkWPBVd3LN8Pnw8FUHiZ2fcdzyQggQ3CHKPxixq78kzUA+lisP0f
KAdm/t3pwXUN5h7b4LMfkNWMObEdGsWIuL9EV+tFgKZtyM4zJ4/NRlfcWZ7CFALPcHvmEg7MgFao
dDFbQFLYBZI5M0BNLXX+Bf8cDIDRpvBYGzJ2CFBSqNpxEH+lz9doJbXWRIjKXtwtMA9nTNrARbkZ
HWfBFtwmZt8CFJrPH8QidcILggCt5l87KNShq24Bro0hxU+BfMCNTZVDGgL15y/0kCa8aUXJ/8DR
bnH20Mqe4FbYPWs3jhLWdgFvX5jPJBXBTo9somPwmTTqP/b99kD3fS6cEiTiTuf9dKrQ2AHUAVPp
xhmm2UwEmHy0erXLTalwCdEe8eQ1JVOO7m6/sMxhHV8jU2iMIyBmagTxS77N7FpyzhdezmNPkck+
iolZglvCzGk/mQlLDt0ZbC90mGfXjHsUTVJrPSnXMQFr3tJfM7Ra765TIGvRekLrgkUf2ljipBpG
kSsEJt2fRpZbbPJyRZCpORyGv77aYv8v3etH0cqrd/w0m/sPiQfX3EIRcmsjKVnpqUCiKjl89/Wo
s6+iCP3rhVOvQ2tkjp3qoG3jR2wNEmwhV4KOd7+8JeQfZ5IoOfK8zLfvcVWo6jV79fPrZ1LzAwCO
M5XPCEUPMiHzVZ5PdWDEPT12orWaduA8SZXnzIKG4fFxiAXMNjJnObc4X78uq6HGUw9pxxk6U1u9
DzowyjpANByvfPPZUdJ0/+sow+INmj0FG46kSoQlSam6Wc02uM7d9+ox41r4HH0y5J8Cv7N+5cdP
r5dqEsrLuS240+C3TI4EiCXm7HeO2pdEgis4IIf3o7UFXa6dVuyPo4rKc7QIL1fEGaa+wFNOFkgQ
xhApacTxkjoE9kyQE/3qUoa6tniJA2xnT8cM8PQL0/KOhn/1D4LV57iRMU7Z1ybe7ogZYa8NdnVf
0IXGiAKXMeycY69t2mA3icf6PmEf0sJ0xbL1nLldW+LWU8VslO3YId9StMlZf+oW3B+n7xbwZGje
nv5U4P9zwiEigmkQCVxo3Fy4+g9IyL+xpbR6RsJc39F5OrmNRYzA8LtoPg8Z9YzrGqwusl2kvkvl
FjYNP9+WQJVHaNFGR+EK9NV5NBQ9n4EKTcg1Nj1jcfIQ1+AWFjpQxGcvLaVYOgZ9YARyi9DcptvP
0Zjx0OIYCK696PaiegSn0zn1FiE/mMkcRakia9sIs87uhv+yUxQppldbi19k6gvkk+KIZFWiwHa8
mwrhWSIaXw39EEiLdPYUTMlckPwrf5goGjQKW/z9OCmJ/yUKj1O6AdXYRQnVnPwH3fv9j6LqlGgL
+EVG1eQsg4HHM1xsI/Dmb+QeebW+Ab8wRlWZnnTbN/73+tayynD86dvP7lxEOQwsm5LO3gq3ccBr
tyH7SaGcNWwjo/lKrsj0HwtM9ABdTqLWGgCI4/PBBaeoLuto/TzmTwyUCHm3+hGLgpdYHsDMz6zt
fPpARVA6eEa4wOtEACqD/t4F2a8D+jh6zsvV7HDnCDtZd9+TnUvgCIexOoym08AdCpR1aRNhSt0o
UlgHAbE1+eHZvF2yEpU5vjFczRg94ogO/nfSbH7d60zO0+xq0v89zMBLg1SwPxU6OoO8XpCgJ/vc
k7LVTl6uwiEljj9iel3u3w6gMM2xE21GHLPraATitU83aToqTLX11Fd4lEwTqnkZ2yItG5ILe2gB
caeCcbgAmgVlEd5Ddm6lnJd93ywTI+MeFr7ugK4wByf5KqcAps/QOfo6hKN8zjeKlCpKrjqbdPgx
cI/dbJCKUG4BNITzSVfgP1Wmvu9gtoxv5/k6gZ7AZdSFRlXmqiR9sOosbBZLSNH5UDwUg+mZADmH
M9qwpwM18FkdiIipnKxe+E8Ayvogk9AYz+fVv/keMwBcCz2I8h2I8HmJEOWFL1/8LMKi5lVbw/HO
DPS3ASlnN9z8VTo1zAdTUaR+KkKUnm0WGUQz+As7rZthZK6AZg1h5R8dPkszTV8/28/vnumg+REV
a7ABr1ugIApU7nENHoVW4l+RGATjTWOjhv7fXWd8oIlbdoUcCOGjPRnLBbyx1Q/dy0CF48Ve9R3B
X9bnHEnNoXZacoYG/y387NU1w90WHg/QKuOs2Y+QPNAL2jmKXEb+YUKICJbx3riveL7SgiQJ9Bqs
3ncj/x8r1az8GCAfkHFlbK8xrPZXWH+mk1TsH0F68ko6RyWmA6eorY0HdPqZXDKDOMjhUAbIxzIf
yh94mw/wNCIc9pjzrZW2KFzck2FSESeg6Mvrr3405R/8s0v0MqkFKJD3RBjOBy9UdWEBcnJGtLrl
U1WD3SIlgbdyeCgdRYv55IHSl/LnAZvq/IfnduN5tUMs40miJJE1kNeuC5UMys3vapHReih7oDfG
vOeN4C2DYWM8TsJ2Wfpb2GfnU4f73dEqbxTyPxLISTvP1vdVBc72y0ZW/JQFT0C3MYuFbfwJyTC5
ot4+7ELPUBSNZmRDMMhdMqAMSffi7oXub4jpoHAzwRW6x7u4IXboSDdhFWjjqsJbmgpti8PnVOJL
rWF8gxc/5QUb/nA+mh+FLOKMIIUTPjV0z5bUKOGg9S6hF6QbjD9Fhwddig/IQE8oCMqIyw4SR3xL
Nl5EgZD1PQtRBA/eYjCnqKd3GzTXfIIODhX8lTU74vvapLFlMHbpEJq513mcyAvrxaeGQ+UOW+1M
YbZRYHwypR6xocbqDH/63XW1y1cHGfXyp0HPLn8LDIXRd+zE/A2UlI2CkWgBDV/VF8xDR15GvYMy
UCvc73HlrcaYsARtDD6irfK15wCTWC6uGp4G/wbgbgF2NsrE2j9fre0lE2fMhekv7EV+7QlD7m0M
oe6KuUay4A83YX7un3gkCcLcry6hDCBEuMgMhsqiNt07ictqnIOeKYU5pAfzOTMqBNwwQd+egMr0
qMlWP3LIsDSiLZEuKLTLvQcd7A3ObneV0Muq2+/O2qDVhZTL0WrFGF7no7o+nPvHLJUIu9I+/8K4
Yd4NC1fm0JwblAtbV8+GA641MeOTFIjqIR6+YqJ/rmhqqiMnwqqQwujQhRD4+ickFTI+OCVJSgW0
IoBrRim9EHEACAJvFoT92ipQpIfHwi7aMmxqR1zMZU+A/mJhn/S3z3EIBXPOfub4VGY2ySoJFwuz
S4E5ACTdQ6RqvyGbMTlg+qj97Fj0p/GdJJWTJkk1Yp113WApBnf5Qi38vxXH4kX7BZP2zXJCyY8c
T8ZiP4DIyTQP09xmfHP8zZU7eo/IGT2priQX7qgiwXb7wuuARoYnJab7IGD/P4XkbAKKngAO2y0Q
Hf5i6uzUNva+DbIm8cYvUzQ/lsrjfDvMzMJHCSVT1QzZac0lZuTZy2d7wtcfTsAklZVI1iXwpc+f
c0YGfFtXYQCB0pVVb93lbrreNaTrIGzwk27fPcZVznpbcDk8DhvOETh7wFCT8K9gfot0aEzR3vuw
v7bSZzCGvoNq2K4rp7u9aGtIJuWgOmxK8yqXPMpTEa5gcDWEX6cq3cIhsht1orwmUMBnRpQQ1bVo
loGQq3wcXql/UuML+CN2jNaQaP/qsRjmFZxZOo/piDQENAyQdi6mw7TeIPD2rAQuopjKnEC80RqE
nJl6vpyyXr104uos5R1Y874+CFk8kiHujsa3AusshHYYG3yMylnKK5xCgiesAT2bqc/R/E1FWLNB
OMO/iY5KDhQ55l+gumqRyJCAD7DKIBj4nhTxe2UPtWvxWHmFRD/Sx8rk36/aCUhoUrTXGFo+TzaB
NVYVk1Z/miu9FzzDGmO29m4scBAexG0J8zo9bhfidTG+WX6Ha4bAssL40zMiZ9Hc8isBC70IiNqZ
fHEBEUdCq0Q+n4g67LWEGF/yv40pHziUolF1qjsSf+aHVQUL2eY0+/YGJm/Jm7b6l3W73z3fFxLu
SdiayzcZbBZZ2QVBe7CYWG5cQRHS8hfkaBAf4G9ZPrG3WkW9eDbwmEZ34nCckuicG9x+DduDsvy5
XWbq/83993u9Ck4weLR5fbOm/MjJ+Mgwsz+WwxLnIde6lDMpurSs+7LljeQNnQU93mvrPS6iRp1A
wSlRCNjDRInmkiJJE5QJBd1ZSSCSLRz/JUhClpVex5p2NEgvH4bsd95MTvd66Al2DvXhR6XkGrl7
l/ug+XlxjppWejyzITouOI9y6HWiaVoCOtpmSyn2yKrLmIGt0OhinhU7WpPkTsNWkU4pb20TOJAl
oCTy/BCV5XvBR20PoLyxJaDlOeObzqFHhm37hdav1cs1vnM45spet1GuZV66VTjJfbg4yNo8UP4r
knKOE/tu/2afhiOfKbgS4/1x4QeQsysp9iFwqCPi/EkFwdPwB6K6sJUdIaNn3QiQeM+cHVTfVOz4
5nGSKW/SUTL5BFqvVKadEJxcQaIgtkZ4REag1Hvm9cpYoJQvg/UAEHKDoJYtHk4/qG3E57qmn7PT
+ZzjXYA70hvQ33KBeoQK248tfDTYdKXT9PKlyADPDfieXgehUNhx7mk9hiYHcqyGTi3wIhFRLnn7
nmrgPhj2QdJBp2HeJu3/Kfm0ifc2tlHh/Iq082Z2ATYXs3EDywjYg0+CfJUzwg/MISHCM3uMp4Ma
B4jyJPK6LsY1evEKowubY8atXZaVAw3xECebFSY0qGMMHB6QMT0BT+/AeNfWrFtsWeyJ/29HNBfm
EyTdou3cbeMA/QWHLMivy1FAysMoKJCnOFw4ctmohIW5nrJtT1WXuJ1hpaO/9+9BEuQyGU/901G6
9uZv9k5pI45Mw7Eq9kNOcbebc6AfXa/BwJZ4Y0h4CWkbur6DyibeVmzlzMT41rUJSmACumWGCyrw
TlY+mJPt6B7SRPOKKcXWM8AIOmBqp0KGcvoF7XtTvrG8VDtDMXT/97Znm5hj1JyTGsxd5t2DWqH8
FD6tpF33Fvnr6rpy2LCB9cbnnYKeEt/Yjxbp/04zor0mEVxb7n/lZUQH1xs+Xpz8f4NApEzP1ENK
N6JJx/TGmnZ6CpnWPOS1Mw5lpJsW+TmmP6ipxWxKd7t4SNdrU4+XHEdV2FKPgPQtRVnyascf4AMb
Hzy8LQGL7ifR9a1DdSu0ovzHphXK4avioq8ktI4e8dyH/Kz9FchLq8IlJ2zSpbIp3geO+E32Qnlu
7eN16vUCIatO/jJFLlwgyfBVoFdwMmoLM1mo9n9KL6HgnuJFvd32LuL3gw9vBxLIsriIK415LWrJ
NmxH8mZpPIgmmPlXuBWNDjxHyrHEjueKMhY0GGyGYexT+JoPgaulC7wsIW0UidFbJs12DeHTH9dv
QaoNaXbLoXE5LqEK5BwcDidmPzdNWoOIJ/apEK7MlMGFJgV5YagMcJj1aVKzOAT4C/qOYOgRRcYF
0Uo1Cmki3ZtFJTdHza3S4ngns9sfE3VItm+GveL2YhZS3zaz2Jrsakycv26GxurnSyQOGqCgLD7j
ekYsf1Y2C3NecIXTP23Sbsv5heqJetweC83KL5mqPv2qOe4glZOxJs2rOUie1VLrRp8GsQuu2lmC
wFuVB3gQjJqUWbSDDS34SSBtPgeLIJkxf9EYmPvxrgSuNqquzjuM/o+fhVmbeaUQM73fFpLORvfg
/Vl1Hkn23GMERwer93pnV7TfFAIZNVzmL7z6y3VsAEBTTt6JrNSL7wt5x5aH2nIgE6f/wPshe/2m
pgIiHqwv5/f/TN07+yPSjOU/iJXCLMXMbzKuDkz9Lfznhyk9bh7hBaT6sqSNyxsNZ6ItFMXGA3WP
+AUD514YCshT+FeMrUY62JD+j6N5rCbax+9T2zvHYY2AKanye8Wph+nsP5r8TZIgJKWQq1czm/gZ
Vve8LEHwR8UTdCGpLCioIXj8GdEZIhSMsWb2ZMWuV+VgM9FBPprG44mQ2Ywl15g2DDO1Te4L+WfN
RvFt5PB8VmDdnRw7sQuEGTzi4ndNsY8FIAGYLjVypjBcuH06ot7/RST9Aw0unk0ATipnUWRx2SYY
80utD5Q2mZxuuuWcxVsgyCfMzCumfx+qiN5XZ9uQmgYuCElofXyxiyI5R8DjEHHkNrs2G2nZvqfK
jjHYZ+7pE8dIVvT9r0ypeZXUsZx6/t/A8o4p/7twqOsduQ7r8KeKDrLlY9Hr4b8o9aSoxY+41Wab
NdP6/wzr5EL0jHYNjZ41pe62kgpgkuFRPIMNWGmX8mXEYlQIC+PutJmMN6M9FwK7ZM73ZgrvJ+nj
BmffruvtCmeheBlJe1McUVj7qnMcnli8THKK3tPMCeSAmqL+WQoZ8SJgW7C/fzKw7gPuW0qRmh0W
TsErVP+yZJH5+4B9pHcgIi9hWscZUUaMkh3lNdYBg28fJO0iHQ4pR9EmH6swJ4ZpXHIC6BC/yUD+
GzrtlGLnJS2rzIdkbCvfgsvTPZ5tVbYOwQsYat3q5TnN+Fu164n4KqukQnWxZyHqlFKqNw+254uy
5ATsXNeJeDGf62IPpPXwy9HVTpzo25pV6zZ1Akaxh9jMKdrBYXmk2RfmeDsJubM18TlPC8R6EVq3
71qBh9UGWo3Z5rGtanjaL+uUg/xJb9HcmkY0Vhy/PYRB6QHUx/LXk5IX2icPD8MJzFz07zh1KATz
TpHlpwiAOwJ9TOzY7FPa1mDPJ8AQSV/2TsUDcy+ksBNaHYCNMavelNiECetsl0HYEB7Kf4+3oWTJ
b6QkQOvmRbGt1jWrlEubM97k3aOUr7nx04xaPJXLEzrtV5exEz5FlTv7zDijWpCOPoZwPjZQwoV8
qAuQasTDMIglpbPvWZArBk/Q4WEqn90pDGE/4+icZUQq6sst9LezXRJQqv/EclFJDUOZxswdep/E
EF5CEENrNdldSVANTIiYamsHAWYjgQ8NTb1YCvK5MbLYdiBxNdNF6vijiO/LDBAL01qUQXWrI6m6
mPbEJN+1JpfkGqiiaycUBOTEiz6OG+Arb1wYTM7t8oz7ATaJAbKwn0e58JfYbx7bZkr+0fjHOUkX
wQ7EFMIcrahDYi9cnUeRJU5NbH1pjLfi5uD/6yjEFfTrc/ub4XuZEEAj/4STDfZqd4hwYDpFfFyZ
I7iygGnvzM7d2GY0sHjBGXhL08oIRq6dtrWlDIC3VOhTnIgkA9aoNHha6qUmODSo/tDW/JX7jRLG
jzYp3Qs86aGDY2Vl6q6EWPLlojrFpoU8xGOq8H9MjDKSOz45wPW68FFH0hANE13tTqLYUKuSeV7l
LHBmiAQqyaRXOb+eW9hssB5I7JabIpdSZyS0v7bqL4X+ErC9/Uc2+W68P7C/c7O5/Q+4n9ApQpug
y7UxMA8mnhD/wJFHT18MjbrJ0y0hxC4aCz837amfXYhIzcd4KZHYxpIuANjElzJvkpi5Bg1b1gzZ
UsqkYIRFqHwR8O+Mqg78Ij8MiWw4ZiQctx+m35vhJyrrntQrCXmb52v3k17ZpDHXkZ1v8MIZmqZf
xiEr62S0UpwUHYe9PcNDxBMfI5xU5xiJLjI3sS3yxWCZ11hLOg+5xpbAszIfaaLOIMa4Ezz0jmow
xRXcJumHoKvGCPsS4591km17yg1eRQ3U2hVH70eUJMFov3DAiVzeg1vQlhbP/YKQnVWkfq+hgR7F
eLs+vLUzV0mb3p2T4Y1f00dTSdnNig90qz/XZcjk47buUeEoAemIjzXEytmPGXBPedS0oQ+twcPE
NegzznKoYM/KMoM9xIAJ89TVuFc2yPdI6QcZGAaRKVRaFK3QKXrIX2rq0gIcBFt0gIas1+pLNd2w
uJesn2EPZ4RGKoNvJCnQvoqmKPmElrv9B3k4kWQLVybYkslVfPlVCrx74oI5ji1x7Ow/WW8BHniY
V+tucN6o4H2LRn03xjrjR+GUqSl8MtkjJwb+a3QDiH9KoIkpW1UKFHYcnN6VgyoBidrJe/ouieT7
I7UOcn0B+hOe547zPr04JcAiNmRgSnmQrk4dcNRmR/RlFxtFNthM48Iq02PCOPqeLqROzk3RDjXS
N+ayQTprTzWKKcTj/7+j4ADMXM4N4doKv/suoawFPvDLPsbLIdFOc2BCR8UbeoPZlyOqfTVp3QzW
UdYsGgMGpsX9IrIYZeUw8w2Ssq5rytSwLd3ykBqyG02p+kWjZ1DKkmuYDBv7+/xLe7OPt5QvR1y8
BWo9qx6gpxp9VGQ2E1CowVHQYXGRJy+vpLxwU/VREHWekBSyUBTlPEoEwWt49ytHoLNERvNWwxu6
lVjeFcBDy+jwh/QvB642dot3UeU3N3trPzAtHNwkEej5UCygAzYj6D6nx4mMSqkc3/kJtrTtwMj6
kwfHTlsu6UuZHWfx5lVG0eU5Zm2SghRx61AZS2r+P0MTeWXFer03QPAZLIVLOzsPBDdcKAjDGaYG
SX1A7qyp3mouoQePxdXd42RkKBm0IrBiNz85V9xSS2+M0y8wt8MsyLqApH3mMx4i2GbeJVvoH+DW
9pUXJbyt/F5fVGzDJ63Bt8LrPxQMr0opjBxo9NvuWxZxH1K+uNuqM6pv3gCpSWOWztVmKczI5X20
KXUT7f+f92SdfCOpuO4Eh6kMFYd+0h2/dDv6I14fKx5GnMQoS11EyYEUuDMqLrCCT55OZphdNp8G
YQGUglLkSFCUVsLDlVFA7XnbEeJqdmJaIVIS6XlOFqfGkzuwiOqZz8QRRtUowCMlN16aiSpBrld7
GWg01aV4K1k9+f0LxWhpugi1C26uDoU2sj4lQniYQwX1BDe4tb/Li5iMSGQxxq3JL1Il9TS72DRr
nHUipGDXbX/zriFHDBacVAtSxjfHBEjY53/dXrf+f385xHt+O45bS+11IkNJcaF5U19xib0UAZtz
yCULtgLQcSOfxtyqVlN/P6PhwdoUW637k0syDDNurLKs7ki/kShdlltjx9MOFtVzzABH45lrZU4C
CfUo/yFP6ddiOZB9ejlwTEqVE58WzaAdaNf2YxiuU+gRpre4Sk8qrQJVPV69CZabi4GyxnQkBoZ2
tU8MJbiloGuwZTt89vmaavivrE+ZnH6S8jQ6U5I80+QVMFajRqnAPJnLV1ZKY+pevHRQYMazInmX
mVZYu/s8nWsPKQ9t9jxpWpjJ0QKswG0diJ0eKd4jWh6NHai/VdKZeHxC6CpLLaaN0LTyLYl7RvTt
CJhsdQ/ZlcxA+RfImWvtRNUQ6ZZHPPK5LAbztL7oqsTv7wiaMMwAITZM20t0FwtXm9hcSHKGYH4T
+oaroPWRa5q90g7LNEm2RvEdp7i1B6+vzDbqUyOcRgc098AEYXjN3S2o2eTP2YArLrD+CSt+SSIT
aBL5tJ+U5n5vCdJURlQUXnJPnJwRBf2qdh1P2MC48I0ggRi9DKfMhBEwr7lObM32hnQHVPH0AeJG
gq3d70PiHxtVU4W47ggPrhFiF+BGmaEYIx22Q2NUnzg2YkDPUYta8ej1frft6UfcTae/yGlLtqJw
4rysHQqd99SetUdmNMwhzAXrPmVT1pPkz4RyenAjOAARtObS0NFvFv9xO2eNZDG0VHC6ijXJSQ1e
QGoUtv+shgu5blYgcmCFkS6atFpAjNzAaDuGX7ltK/xXnrk0PC5rBy3ah3lXPl6zCdCSSburWIra
/6dGrzhwdefG056ZmnTCkKBseTEoc242RGWI5z7WJVy22tzwOopWoFYW7/ArlWkV6uXuth1wAlPQ
CL8qp1OWkDtI4cDhT9jyoclWlSW/3qjYma1fb9ECZnAPze294cfeuhL8G70mIwPfuVQ2TbelIqNE
INIcKh2V0F5d+8Pax8Px6WHm+xU5Lq2sZ3yT5YEyfYiioR0g9/f/rz2g96L4EGWYlvmk7jPD/433
09srsMzfDNiIUDwWXNTf5SU8K3BgvxBF6pNn2mXtZLv9/s5rIoFbO1ON/ZiRNcYL7zXR63aoPIHp
Yt626GiO1f/HNJVuu0TXU2+1dkG+OEKy8rhxhA0QzzXGnUsEpbJIFdqPyvyBzuqIXnn1EqT6hEee
WBLRBXoLXZjApMJF4O3vesy4QOUGeVeFTbAtyD2Nnd+12jTmEjPRRcULfS1NXEq21rX/LsHHf2GG
VthU+ouwhZIZlc6p8ZwR5r3ZgauEYhP5m9ZJKKhhGqMACKcCCUhZFFNlCIiM+PNcxvl4C1W6n96P
NAWTR3yhwnCkkoiM8Fm6j6h7wJMbANG+2QO2tTUeVtAb5HR7lArA8IQ2egZdBgZ7saQT8yS2bSMU
C8/qlEfWTVY37O+JafDVhNdMBHH7IHe/rMf2+OXfcMNp0VP3eEXyoDbbhj3niPu+V57+HWOlYZ8r
32/XlkApPLlnCuB+SlAZ5FtlaKT3RBH7gUfGM8WSd3w0nXtTqeOPO3mt8qWVGeODC6554zYXE41z
YFwoL6U+DlsYwfqYdtZuHbYXbm02OuoOGnBhtw7wTNxOSdLmOEURgds315g0CR6ve9ne/2jFLBX8
KpGglCRY4z4QGx+tAOO9fYQ2xXejFLSavmFBfR4JTMcITQqhEap1UEJXpjTb6M43f6p+Js0XJBfk
xHBCl5f1dD89yCVciVyoo2mZ/HlicLbm32WiQPgoUS6RzDXqqRrp7lrk9hllNPXEYYXYprnRV2uo
xls6aHNBWHS5fyhV8a0k5uxdHikY6meTC9RYtzDJD6mBrvxCq8I/2h8z7biGZ3UgE/c84aooTbfZ
Jzo2EwMRcBBvidzyRaYILpNYSCpXyDPDpUYBjJFYUNuGp792fXFz1CO7QO833ghrJ5NTI+h4ZF7v
lDZnrgVnAFczX2NCo2qtRk3TCfuOG0u39SZEzWc6Ci7/fiWcFoUorimhR7bcdzTQO+UwvIvtsRW5
nnIc8hp8N7ZZfhgUInOpbkCqaBijhKwlf1P3FHwaCMjSD7NJSjxThwGAGgxDfIiOybcC5LM9VnXo
bJJ0jPu/uu3/bfCesXlcSt5F5+7TkpMvkPEe/2GoJ3btKRzuGWkzhLiKvdEZKgGHRJ98uOPRAdus
8uWKPuUPTUaq7PBOUXXTCcCUBTEckvU5wLedzpxdJUZMbPMW+bU0o/oGYjdJGAtrV7i2knb2X/jE
x4kVWE0HG+vaWRwlMzW24yyty2IJXx9Mk2dNA4UVsD5OcWF12ngIGzcBgyKGczuxxkcJ28KXvM1T
E5zBN3OtKDp4D33jVdQ3+S33RCZCiPHFzhXYYpulxmK1jOaBd34e76vgz6zzCoINy2uD3J7MT/8u
BNe3ApT603EKJSEOrrvlbmuOEaDndQJsK7nwlrZoXF2+pgmhkmzSs8g4iOvtqN3oH4nhkUg8rR9V
O2SVBsRXb8IEZfX6pvkuirhwsRcXPFGf+gjsPOIezzZsXlFkEWSqKmAB3aJKX1G8zE9FgKZY/uLU
RnlkA199MxK2YDfNdVnF3t49nnRSenxWJZcaORdDV1k6rHXwTsnUhLI2oUFle6h/sXX16iw7D3zf
uHYAASG4jqvaHXm/de12LtgBODKxAnjekwjA+D8pIWfXcX+OZLeJrk+NND57OaBoruRAHs/zMO4Q
3EjO+/c46jfFyFRUOxCDAkZn0y+MnhY8yfuNJ+5AgRxpajfwzJNretli/GOdPGtj4XvyZ1ikzURx
PwSZr1Wzub1FXxRDsDctLDmp5mKRHWGgLBkoJ9WE5e/jfHv5KRegUyOnePYqGb3mWk8gp9URQM8E
qq/eYbIjYxEc27aFdrWmQ+WKZrs9j/PybSCd44qkmN4DlVRmQo2hrd3BpgSeXgdM/Q125PesSPCe
XMH4pfLdyEdsK9ZNQvTGugFJiS/xDT2zaX9Y542LmLGsyaMsGa+qwbIG71wZRndm+HS6HGGbrvdh
frSK+HYuqo5mS8e2Pb5RGbFMJ2rXpdZ2REAZatSX0AIwXK/kcHG0CXjdxKBZ1R4uMnO/GLoz0uXw
9uPJ+51PyCPjDbcFs72yJ2x9xVPpqyBnKsCVh8+wjA/NTL3x5Y7IoMRTNtR7yjRlUvGcow0L9gdy
BN8fxHN9FxZqNLRpBeHZ5x6rIjkOdfLIluEkMOyHqYQ4SbPV7AGnm8b6xySyQ36vRggi5Y1KB1Rv
TKo89sFmTQyHP/g3oMcYHLNBDlYHBAOg/2NFwDfyRqHwwpVAQktN0oV8gjQdpKzyJ6mmdj7TOcsf
8/lZFz4++Z9Ag0A0S7xvbKN/b93as9323eKnQWPLgs6U4455oovQz+JY79BY8fmCf6PwOsl5er63
+4ZMP/sIxmWPGWw/6/hKkzy3a8k3pIP4xrWS8pZl2Ew+Ctyp11GbEeonk8O9J0W+3cns7b8Yr0dX
4GPVCgIjCO/ST/es9Gc/g8dBB/pGa6Szq4Z5LgaoX6pGaWlBBuh8b4bWgwaBZ5btmuicZrtWsxKJ
IqPwYywv4kb8rt3a/GoMObXP79LTj8/nZHVfEQ+BpL/CWyTaHRuzWAv57zquLSj1rOt2edxskK0B
MaaVC07siSv+GGkuqslSRAMrktZrv31FrNRoIZZPo4Xt8DWmv6IXzbqcJHd2c6uSLQYjzdh9D755
ST0yU/RnlVEauUXPz8DjKcqnvo4crktcnHh8VCb/jc2fHk1fv7LWWNjEme95go/Gk1iSYpWPoaPt
UbDH6B8/471/I2suvqIhWTHECtNaN34dcOWwY9+Nkj46tItGwjrLoA6sddVrpyJ6e89c+MjQA+EE
5LTi1MrQzRlZysbHk0H0xGix6YjN6i9zq255McqgUt03C4ZoSaQV7RwVSu1U9xsJcjNAYvP7XGbr
OF8qbfRH1HrpXYSEYDuBCcaIssRxxYatIuSIxnIk4yomZBgXL6Z2YsFKUhnGNtnuJB90eVoj8RMg
HzQKdWcVCvLsSsLg4vBhxXFx4NFZEoBbzEYcBx6vDCL2+TDDChPz9SSHLL2evrjUANNOixlFx6ne
DndJDVL5kJi8o0usZBb9tr9lX5Dp17Hu9FKT9D3R83xJ7NKhfERQXyo3B1DRCEiUUc/VSTKUp6uR
UbQ6pddfKWCNnjU6H/+VKGxQs+iTaCXfnUZpJ4obuLiJWzF51dDs0Su1zEht+8c3y/BUfpL7rBH/
2unN0njRuf3YbfvTgD1hjT6Ze+7oGVsEyEMILtqvet2w0cxT9tduL0se9yoUpVWLeNHZANRoHwjG
JPYp1N6nLJ5LjwUb5myEU8cOEwF44BVssowei4wC9setaLle2V6Qe3aEKt39UB93b82BQAi8TVCW
tCawMLVz+ZKCQq4acfdn1ydF2l5js8fdC+mxgpyJh4U5DvnlR6lcJW0XLNNqSbRxXgkQsbUCrJXn
FUKusMgWfvDJdC0OVU2rsCil9GdzuK3WDZ4/p0PjzrlDLMy5eI08zPZW6joTSqA4IyUyqU6UNo9F
5lvD2YwiDeGHsGwLYnc1ESskTimdZqhdlrOwwW9KGZi+7Jl/8YjdDXX6qt8GPUu7My1O131dnAt/
Tl6PRf0m1s+oIK1K1JlU3xS31t5YhETlaDR3uQCl3EkrL1Yhn0PGHz8yfCGyGOsYIuFCHjYCYcN0
SjKg2zMmZVEsVBksquPlCnJtAtkC+4gPPDwAVND9EcIOwlDtoLT796P26qbJi4QhsBIL9rYUVesU
iTufcBKviFXkVfsfVqgNL9CGH+RfMRZ2/oCnn8IwYO6L5/5awMJD+4Fy3ZDXyOMf9EndBkRpTggK
cQZdKjTRD+nyI/zQtU9eMzijWeiGlUFoM6zdaFVaOKfVU7N6rfPZtdwqY7LLLLlOc+JWu/15apOi
YRgA78gjfbGjZ5rYsYtT/0HF5/bRzqHOF7WrRUMA20oorfwqGqyWqZVi/tm4GR3oRoLoxi6sFGfc
w6Kx+tfo6bYpdXrY6LiMBhpavamQbteYpWR0s0laX6dU/t/K3lyAD+nRRV6I9a39Psizya2kITw3
51z9pIEXkV9ZQGhawZvash0YXrVJK6mwjG9MUGH2kMTlfmXTNYbW+Ig3kSL7IhxCHmJVb/1PCKm2
4Yl1Gyxf+HW6q1GdRZClbHmTUhdgTBDoHALUroc0YJ6W8awsXPIXc8DwJjWFqCK0J0aQc6IOyB7l
bqHkzZphzvIOy/mBAbxFhY9ynjhVYNBMpHr6Aa5cfGUUOTbwlpz4+83icZurHt/L/XN9HYHjE+/0
QrKgC9vzJKBCbTigyzkOaipvc9M9DeYwsXobnHnLUIHOyu5BI/VQ9x9R2DlMPQdJb40NB494paFD
IdAbhBeKxy/rKqnRRaL5WaPNJGefF8Xe6qxBZc0FsAHJ06oB06cmqjimN0UjTVKgaOvDIKmbI8NS
Yb+dSX1QZDFmir5RiP23unxGlN3FwZWI/BIF2TPsS5W51n8RW55dUcHDrUKZyRW8efX4FBn/qDJk
MsAEsiZ1j3Il8Qeumy5Hzh74AVTvzadQmC99/fZHNYxHPGeDBL1PmYSAX5fYi0Qera3x1gzIhm1a
ur8/fuVefUfU9RkhVgtNl0reyjreKJtK45BvDgVD+ewt7/fQNbokjwbTc8Xc2mHYq7bOgK976+ng
+c057KibUXGygaKV5JjXCgQLH+PywDxXHjghmVqLTBQjXbaXMw2pgvsvUndR5CprdGYqVLarZL3j
rd33KTetLwlr3Y+Sx7tMH1HGoLQg+mgIGgfu+QEvQTLs5PJx25tSa+X8JRnwgXE7S8EeZ+c2TWxW
UA5eFvbkFnteu/Wg8hrnN93URchKW0Sn9/WQTapUp12GbSn46w23jS0rPlPSt9njDs5iWBS349B4
MmD3/fyyjWRytopTSYIkBzqM/tnwAcikXma4UKcQoIMyM5NGib65QMUDuM52VKjyftr59o6Lc4zU
SoORJSYHsFpm3ZzEjxWXwQBRj3RdHjbj6NdgQzmrZgqsR4A9CTLLd6FTKkBi4SehGYGXmCIDRNUv
HVmf603dHJ7GGR7Onxk37JMGIFUCUJKlO/CQhFvPO7UfIAeJmOKWRdtQJz8JM173AwqFckFVRPoG
g6DmbSVgYam5gAMMtmH0BJj0sD39G7WNMaCMKn621lFMXcMZxlYtJweLWhTMVGD2OBIB4x1QR4W5
c2lwUOlZkQcZ6HgXpT89YL4G8u0RoaJwl40zVM3zNr/1OJ75B9afi2C1xe3r8RQ6gzzEgmACRcYQ
SP5MzEmvQkfnbt2SYPjHEZ8W0ibfPjhG4/QjNO9ocBPO397OucS2WKuBUCotdBZYIuqrmrhjuGzu
vDQxRPSez/vd48HHJJuogzNSZJnbZkyX7QuccBm+uIy8KG9W+H6iCaoEJdiwRIu5a8A9yyr7dFE9
AVs9XCfKqudAgXhnimWB7xwhH4eeKCANZIsdR5VbBqWwFDlMO1R8LLzd2KmDJJkA1xcgNMnLvG2F
+kjEpxBUwJazbfZPzqDdwdNiogchhOEyVngsssVk0g8POMa/xN5jq02GnAFJXJQ0hsD9yHyPRsB8
Lctu65ElhaNhRjGwSTmzhqE7l7djmEWVytlgk9Vl19e95Vu7kNQSQfcZbzKxwVOxA3BmmdtJ3yO6
eRHwwevItuNHkJlR+cHA/xPBP9YINlBTpmCH+REtKFcpsT61Hp4rSsLxoDtUdjsBI1mVgwqwp7ZQ
QfFDc/P6KImTQzf+dxRKu/IGLAJE8/rLF68kVdI3yf9Q8EDotn5OvOrhKmd6HZewdAsP5RgXJlqq
stG/Ej1gK6M2Viqd+uZVJXzsiwEBg7xc2BglSde+v7mxiCInMqXVUjUEDjVzensERlXT8qsAgkeC
2mgYklWL4vcqZYBZ+HyWdGaqwyEg9IGmk19nUhO3N/avwX4gkZeezykoJUChGG6+fdYjXP85My5h
MJQhTg7Fr/Df+JCBdkGTSqhQbIS5if1VHrFJQ9YG7G6W5cEawfH5pn4x9yYx9piLInxUdz2DQ4YQ
AIW79ju2SRsz9K91U4S9omuOJnrGI10bpT1y+193AkdaGi68+6uhxP1LAbzvKuPcxgtiqggu95/K
1aUDwjtVnG5vcvrY7AeKQCm1+DKJxfwQR75F0c9WRgv//wHfqwMA1+/1/XAO+vBTpYeXPT6rvXCz
TSj2oTnkLoZJnLAH/ykssm5eOcSuIJkTqdT/+Q0ggwQDj4eIWfnHmh1yCHDxMscJZKwh/PMeVDPO
44k5/GCjWnDIk9l9MlYEZgXqRfAop/gc+ygOtA4u1Amih73LR0jHZyg1ayOZa8/yBWrtQfs4+ZWT
X9Zb2iA5ySWpDclRmP5LNNVQmVKjSuy4wGBIwxSKsfCNeMlvzntWGLf6LzfORNvm4aqdxjUJFsJM
mmTIpCcb0HUv3G0pQ9cjKJ3rsjqmJXikG5COqqWDo7KlHlWsohPKQXmwmZwZvpNrWiD1AogbNtTv
buxXmSYCxXygA9xwo3Ss60vKZZ4VLDE8Uu5USMAekXbqP3gk+Wv95bJzwsNV50dnLqwiAdg5XMUS
uGzlxdlWH1Y8SXG5eHKPfo9PCR/A1ahsmCrrlGxDiOs7e8J5LEWcNpU6oAY3HdoMtVNkxWF33NEs
Yqf+3KT/hbFPoVJbjq9CYwKccinipZirTfIj+HDX4lSxzUogG1kjUoriOb+79JDPhaa1xtbIHbCa
sLd62J5UQo60AhwQjgb7WhIgzKXKmsWpCgitrfzYlbtp+2wOlQpal84j7s4OuG3s6F24FgO4sITs
yMXXBNfGSuyQCqsKMvdgBmuFgZkS6oe7ECtxmPUcI9gOQSehJaVnUpAXhNlJAb+gvQqEmRLW7mB3
Y/boqaWLSENYVC0nG1dMLMfOllbSu7tw2KlvX3XeM5jmAXbn/mPl6eRmCYeVAfyPx7FTU0o0MWA3
DxmPaW0TeQOqA+4J5HozVYpbHMGgxd/gpb5vWeHKutvcecc5OMGrbjOumHn66zn9xZTeoaNn/sjZ
ayjOS1INQURINpcLkAPBhwrqXuWO/GsApXqT24nQIw9ORopbpQT+qSXNY5cQwZePugOYV9+XZU7F
qp0C+gACacp+cFPUp3gqXRq/v6xRfj/QriiA+00FwpiKkUxNf1OQOGB5PPkFwMLMZAuOhVTrHEmW
o0kGeXCUyYMbzglV0VgK3g4RpAtvHBUp6156xuDuOO9m0RXxFrk3AxhVQ73J6S8K4rX/gs642Hyg
TWyTQ6fkKZbX9wNE3ruLijfP9CSXw4f8y3ADd8i2e3SwSEAgKN9XC5p0eaqhYz3NxbFXD1z12IbT
wYzu4WlH84TeUUbNmmi4YS6W6wPWyC0fIoAcoqdU17tbYYzPxcAOYOGJR6GU3k7mLoKhoUJWqne1
RpSJSiILMxthi4s0ogmuiBvi1ZiR3hRJBOAPQUit8ShUV73dnX2B8U92bN/2DJNyqYtqZfkA7+pu
CNaDgg9hbR/GEOsoclyszc0qMr0ziyPDwrex1VfyyBfKxXaYkdu8bRpfQAEjy/wWkduQsPzxhB2i
MwaaA+8XT+R0Ln6IA28WZYAg5cgDxAP0uqZ9y/iI/4d2wGHw/TzcUbGAp4gzx7FO/b5NVEqTqw2G
nt45EMcQpKuaUthGZsnQWQAUeUJXbnFsJgBUD2Aq8xaL/wt9mW0ll+E15Pj721x48jh6Ec+tXO0p
Fdpl6oViNiU0s/493f+AanIjJqrcITTB+IV0vUNysw07yTsk6foAUTAsdALSIFZTzoyCCyXBBVcv
VvfS8UFDw7aoFsNMXkbfuszy21pNOibTTb+MYWPki6+YvTlR+A8ImjX8Dva/acCj2me5hTUqJnLY
YiS1TRjIdIZvovAKidSyPGMHiNS7NbbfmRy+yPoMACQvbwMf/nXC8ezI5op73mMBI4x+e7QkAG0x
xV1HLifKbT32iycXu1T+V5QwvjqNJJuBzVbEPjrZnfHZWNrXYS1LLFvaWZflq/qMSQcsc2jC+34w
poTpIFF9ZFbbyEo7XfUuBMjCx9tuTtdV/4SIQ9KH77H6z7p6sCPxIT/Mx1kR3bUCjWu5w3hoBgxm
dnf5PG/2pRAZRO/weJMEBxkLlXRaDooYU7vxgMkOHX7WKpM6ALCJ84grCbCO2JY+sXaMoa6xpVQW
MDTK2UXXbITagne9nYTxnLQ9kCzgGFg8aMYBSPuEh2IYu4w1MysNaT46nmPScsrjbTBzaZAJGREV
58n9NJ3iloz2TEmwdu6hXbC772nwSyAQld6dhYQEnaTBScIrw0X+pcDMjL6VsjNcKZpIqlDOvpIV
RgEIUTxjCpTuWx/r2rZcBr9Re3G6WWeOYeNOAeGMHuP6VvD0/6ej74nINRNkYaird4/HexJQ9C9J
wiSW5nXIHTtygHhLQf9GF6YTeTqCOwbrN0dnr5kVzt0a0NpftO3F9TU5fu1YBNpXudC+NyOpC5iy
p7rM2gcHPLqHP6nP6HI41fJF9JbOpkGD3aPkYygH+GFTXpQw2vX1+54zb1pc5OiDPUTC/cwukjh2
BnhjqzM4guodvm258XTmYc06bPk4JOjvVBXFymUfWRaoYCjT67tDKwecPNXqNGuF7VTZrvuux009
uqXuGo4E1m2pDCstn+I9TtZuQgg6HurylSCgwLKgHtw1aCBrsSxUtb1d6MsBKQ3yZqcosTWfQi2Y
VJ4nW3c1Jqp5jmPu69vW/un1eEScn4W8oon3R7aneleMuvDBKolSRQFTC2kRp/nQeJLBftTZ6jyO
shcrBwLEwxkRjawToDIaVYyC2q0M12DyeAKlgE54qZqUZQP0nC5nVdi4fzu5YJ1N9haNVmjREDke
VyXxtzCOURrgtLbu6buVZ05v10B9gLPQYZTGa4ji55YAtUCqcwDhjIwOOhruZPIaBspKmQE5XOde
EKh3yPlVeAbfGkiu8JgdRQYcsaU5WggQARdqDHXxTxohU2ueBce7DrBk3jZKYuXHkPYzZ6jPmlZy
CusGs4SwEr2pjnq5S9tluUbeX+4y9odTcsvVLv/rPshl0hhoPPvzYxBljhDduvKTw35de5TLMysi
d+Z8LhBjUMdHEqqWpLJAwLXI5nasQK96Wg3hPwREqLQWtAWzG2FiNCUYFYP7853c5FjjvyCGbjcE
bK/x7Vhu8RosUiC9ESDdw1dQpV48adBS+Yw0g3I1R1Y/xljBQBH8YTu1FLuiWaGV39JcfLEaZ8SI
+NynV+2PSuh+44XDco6m/7YaOGsU8vPwrjahoAb2sP35zyEFjzoYD1do46ecWqIckiuSE/KXL1ah
oACkUyaYK2hmW2/CJmFG9snAtVkc0GMyCiwHtgxtUlQGx9GxiKElyxG2Ssq7BBq8O2gp6Wd4Cdwc
SvmKWTG43aIpfSPbJAgy1A/ExKFS5TS8mSdcsjQLElXoLuWHbkwIb+jnfPb/hIID5qCsXNvXVDcj
57ibWNQAKb3El1ZxlaKI4vmrsu/Y2tRfxIEX1aKM6BgeAzOgPp+FAv4+iQ4DzhwWK9IZoQwXFDid
0UNSzwZBxQ4zIE68EwWoGJlgl0SiNiEq1BVhBhKLl3VNjqyvxfCe3KMX8ma0ReAgNwGxqIved8Na
/HjkycuWf3iohvC1sEAAx+rgFmKKXaHGZ4vEgGoY3AacrZno4qSmV4OsjSOsmquVEH2Eztp8lUvt
3f7SkZ67d1tWEfrwEUdqLpnotlWw9r86aDhCJOH2EbQRb1/Xeiu5Kx47TiDOO/iaWgYZy/MUNhOV
eLGeP0nwRZoHEGL+Sn23QHmS/dBaeRQxMXB2k0D6HlPIhQCw2xXqxx+/TwNrLo7iKEoEbqE/ywce
McXJFlWMF9HTssD9CBEb6PepvGGBM4qLx5QG7VGaidwyPTphn43zHaas2cBEwD/T0+31JhYyXr/Z
7d1YLNh4H4vWAJ4nhS6UWdDt3cgzzAHnAY8hng+yuLHy9qAYc/xF0xyDUTAYiMHOfvgHKUyPXHcE
fRdX2L4Erj6pcd0wrhZoLEsKtY9u/p1/b1koxRpfXDPWVrmjNcBb54tfcNszJyLgyQGoGoY18f1V
2/1q4av1TaL5B2RTQ7KMa35TGtbeJBPjCLrPcboF+Vf802s7WxY7DNvRxOHfri3Jcl4w2GvbhTjS
y93tJ93S7j2/Vkgcea58/a+KrEX2wRN0cKfyL1PXA97kU8INf9WqXVAoH93R3LoItkSGq1uw3JJR
g5Y/sO3AW+PC1rI1KzZB3pjeYiPh+Cv/TNkfEarQX6pGWqo3ApEkKHjcly7ocGXOKOWcaktrA3zg
s/Cjy5S2jBwgi+vr7Mdap3iz5khAJk+jcX3+31q8zJjAls9CFZdoQ11Ymhh4dO8dPp7FMxwge6RO
dZm0peDIuA+wYv8rWjXapELIgKDtGcXMjBqgnyflPEZhLAZuq9yIeHqTe6uSRLCDBGVDhoBkYI6D
XrttCQWCdTP4W2S7jEMRB8+HIlfj+R1UdQCTh9RXL9rXiREbGpmYoqhvM+sT5qaO+4JqAXeyzfW+
qIAA0WnPepVwiQDnnOGT1uLEwQrQxxV+83PBfYsx5xDQOgIq/M6N98NKOVjt77RJ5Vwj5pwhN9GK
VpMbx5Eot9bFpRwTLnQB6M8a5XPmfPOQf7Ob20tw/KwmMwxj5A0w3N405uTnAN8Ay/S7Ao0gHTxB
WiP80Ocv+7VdN+1HqhhtrOnbt8UNpIbV+312SNuFYFEnjS+fTnz+jMz6JT+F/mYMCBgf8IukLQDe
Cv4Ua5P6v2EoxeCRbVlgIrRhaEQhGqxzbYlqmy4Efj+Xu9IhCOCcDUU8vVrKn3XCUTQTzCjE8ILt
qNetB0ymMJxdZNBvJJa/bWFvN1miyfyi+6SYb4S3leh9MJ0Z8Rlt6iXEZI/3/LN02Dz/ulW6UI13
nTnTT2/fKqyR2IRWAeJHcFCNFCvpTjyfr9Dn4545S/4XlVbmcTP8PWKXZoG6iZclY7kTT6pet5+C
7y5ImlwFWtRIyMF3wBNKDS/Ah5ivSMmna+nXqYdbObqW5+pZkMalOD4wdcdrBmPmXo+2qNIIBkEL
37cPu0VoHlC5eP+QejDirzwHJT53+GfzWriN2g0lcpUzzeudQ+z3TaBxEf3CGNByxjfNNmNzm8i1
i9vW1Fg0+g4zBbY663kDIBjNtAi924T9xrzNGaYhN3/WtKKW4IUVbZqChLuCbtHVpf1MunozV8MZ
gmJEK0CvvsnRDzIsGr/EV+wXOWNiD+J8p8FMynjKMYOqEy20w0ilwNvJijNSlMIJoBzRFV/I6WJt
RwjN4Xzgkh7Xa37JdKHO4i4be4+KL47Uv5V0xG17pw7o0saX2Ha2WNwHWmcN9FtC3BUillU0ftdZ
2cl+4C0BU4/tEyem2uI38d1WzNNNB4MG52KUnThfiis7NmxrQDQM5q/iOLVvX8BkKt1tF+oAaR6F
6A8qDioG/nzEXt9SUu6m6hghVsDD21BCcP1rUfbSToBrSCeiPh141FM2rof3K9b4Uxo6ieO0TFWU
1HlZuOBh+JCXsL4j6f4s2aZqVlhbE7g0HL7lO3K2+exoCNZUy9OcVmKH1U8OTq4BBqdnu8IBs4sH
hTBTYUBz8DJs3XVzMbRpNK1P0MWmGiqYn/P4fyMuJGOUQQvat+bioBohIW+9+nXYBJDEzq+z09ym
p+3rRYfcqO/Qxg4H3ng5q6pzwXrZdde2a7wizXkWkuzvBlXkm6ZKMrwpOAnqWJ3atEwDiiw4w1En
K8/fVSIFjQ1LkOA4GGorq0Z2JTInZr5psJlV7le5+KUwyYg9AMAjn7q97msnFc6o/WL9q55PClYu
Ar6Pt0FlL0mENQYq17QfwXnlXov1IprHQ6ULU1HCr2jWpVBDJb3GzHGFanHLjbroJGHN96psih96
SHGf3IwTW5joNTxduh24G1zk2UlZCMgR+nmeyRiX03AqdujZgwZ/x+tWvU6HH8lJEYKgOie5Mm+l
sJPgK1LwSw67EeFzBuCiE8XiEXLzWXJy6sOtl+nP4MwqksDJUl2cqP3vJwsnX/Jlc+ek3K8Sfamd
xYA2mNRDtJgZSsEfmxgKVj1Q23tYg6nCV/y+VlSMmktJf3zNBJRSsVRELpvC+bU4cPbUeLRVPNII
IvxOR/TqV7ng5kSKOvgvsa4XDs9PS/s+UiuYn8kSDWoillPtoWN53i++9dcsLg/a/zCAQoAK6WjS
dFoGrCXj4RYtflEIBMTjQptkrPJ65aWCISCpPf1ukiZm1eDCTHsoQ8CYKBI6UjASFtWQAk+YIOyR
ff7wW2sdizYm02EBnSzoR7lByYR6NCVPFlWbtYAT0HDWZUI7Gwpk+4NnbtcG8Sb2ZAw6gQxCtXfE
DS9TbsgX/BqIvYsSAfNZ/RkAukVekboDFsp5kHSAt4hq6nuh4VR8u1KD4uPWliRjVvv9tIFwQCK4
pBnfNwO35lMVWcs1DbJ1yCgZKzg/zi04YHIyFoj2I2n9XxtgHOyyoryQX4SuX5pfkJa/fBg3E6Z/
0O+IiA+F+dTyctJqQxcTzVKEejMPeecf+XFT1a6pqAu5gRl0ShUaTeVeM05pgxLny2XIR+GDOAxI
HDXjv1m+xG+qjRZ3NOl7n5+swRL3XTq05/oxCHW5Cr3RrDRfBMoAwI7Rj/Q4V+5VN3uYD1NQ4Vqp
tfO/6yVTT8I0d7yQvpZTzMb5Nm9wuUXiJMV7G4Jmb35LmNi4rytgzMac16fGrR/jdiKR3FX6E7FJ
+gCmJPXREpj6e9s2UZTpbllo5d1AHZcuGDtVHHmr6xMg6xwM8qsHuBiPwpfeLOhCXpay/higYhoU
+1uJ6VVZreCu3F45zgsvHTpj4xjh2ekzbcG3iTeMig3YivTSr49IwF4BhQWN10iETaMzBYnRMwBD
SrUoCw60PnNdqVY17yOLZ/VubSkUo2Wk40DOXKnvF8HfQ+8eU/e2VqyDlnabhmaZo8vtyoimQrzQ
8zVvIzjY6KTLWQP3j5+No248tGGTe9TRUWYf37ERyPnK7KHkhaffQsN5AQeod15C8c5DxlMmmi5x
89CMK70tR7jZZranwNMW8+TMVi1UthSQYj44bal4L9cPFLy9kowur0RZE0yQju5P9jeuxz7DrAZi
lJ32tZxkQekrMLceNSMsokefvAYTeqQ962Mzaf4lMg7vn/i1v7CuD3wUNrj9cHBMZmRhCZpzG7Z8
CZE0xtG56RRVi9T3htyIDUd4GSzOjQuS0HHL34l1HTQAmZGmgKsEXIT/d8NtMnTSWWK7d9T+brRZ
6bc+c9YTKEttuchB3AFEYoiiLRU0Qyn1SDXJ04FnPhmXCstmKecAXtyzqoE27Lyi8d1k6L3XMIfB
3cmHoKMQdnlyKQplrOKKfvPT2c1matrw1BYThRQs6TCnx+QP0fg202pL1tGlMm7GH/WUjhMYI7D8
KwjbkBHkTdMIOJbcGqoerrNp7fndjli6vtYTqGekXUxjdUJ2tedTaTBK0EqEqXQUAvUyToQSA+b/
EVnQgFjlBB8zG3SgPJGUmgnXzI7W8PZOUkKHxdf0bkiqtUx1uvh+woJfQ65mR900QnuPPWxGdBMf
Drc5ur75Nd3Wh8gKmYN3lYqrGVnIUdtfhFDx1wtoFt7A4JN2gmpTv8WV9QFCuC6fAmcPbFXNIqn9
CzSPMnzCCB8HTlkkVEM1bmBK8gzxfPjKx1AnGDiZDhcyNQzX0CEFVn4nMYZ0Dj/Wqg5djYG7nrAP
xlwUsvioDLPlUfxDlvbPepGIrxQeGRG00k0hwBjJ+6T1K66QZ7XeAjXOShXK7IsYyC6WHBipYn9d
GPhzcbRVnLF8Srbx2QAIxkX+me33dm0alSQlheSjTp0JobiMAzfZeC4X9aH2fsWwRgEqsRhCbfPf
5554pKMB1Kw6RmNu++TAZ26fUrqpmCZMi+pLXGAS2AQIh9o3cxfneg/715UQ1Nls4umEus7Bgvyf
8ZnrqF+XQYTbbU0Q7Nd3/qbbCZrKZA8pZOzte8xKfDDWGS1xTScwghkGyP4SMU5hB9YWhYsEtgwg
gmlg8K26oz0M4UDn/rocoPIB13jO0WgTA/lPc1LL5jriCgAIrWvOfhd6Nh8cAAe28EcoLjTDvC11
qBPZ39SFLhgeOkxggUiaBqhVF+LMht0I8M+x/ZKNGEW9J6YF9ycaUaM2pGUSCcviO71aIJnS8wZk
o4jHa8heKq7ODFpBoDWT3D2XzCijEldTWg7o2ROLk/aJN9ziS4EswJhglKbn15fyLVRJQwlWEad5
YtI0EvbRPrTZannpxgIZBne/VsYdVYBWp0Pr/xTFB8tqMBQw80jNtsiEeWxKuABgapXt1tBVFS1f
fe+elNE1eRPNbyQJlt2JH0BE+3A0ARLPH2fCObg3O1YVDEIxinMdPibv0QVsId8LASvuC4abzrC9
l95ntkpMMJi4iCfOCggL3l0jxsXbqdV87pRAvmoAJHaJ1MgfGNZtW3ZGz0CZkMsg1ikisqwGIsVH
VwdGxYr4r1NIf6RUVXyncdoiEgHBB3H6xrN4C0ljin6ML4L8sqZM+1SwnImLp6PK33llpgrg5GLH
LX62xkd3KtkACfVLUUA1TOdWj+IHqCxqK3SesK+2Grrx6O/eWepqUukJVtJoAd41+kEmsi+kbC0U
vvaqhN6qt5W2NDAq5On3DTVWwUTMTWQ0Q/P/C680enmvOngBgWwv131MSJi+jgdIZB82tpTUYiZf
b8oM/c1gBPmcR+Hr6TcW2UJBfG2Bqraa5x+h25KjabWRFPbKUl8JnQkUh9RsLSKoqReOwf24zM+k
1/EDh09cYNdhBvZqS8FUZRNCP1cUAw9ea+NiEqyFs1sB7J06SU6S6LnXP7BQdfkeE4Z6ad88Ff7E
qjREGKPEWx9wgZCzI0gsNb9v2Kk/8hhl3mHv9NllQX5i0XaYrHh/qZLF/PE91EcaRut5DbyKNKcy
/yN06QBFw4/Pns5eFok77OY3MEylGN1LQlcjL7MyxIjCXVHzZ8UXRlujD0XLryXQg7SZsO/TMHYl
LgL31LNXjdrafRdb0MCHetqTp1MrdFRm4/JrWM+1wKpeFta6/l70SNaGsTmi6kJQUzec60xgZIuQ
G8yRgdF+wyALmgI4bMHNR5YHsVLv97SEAjKE67XNdHrNXmDIltzaqpkpvRYv+3PZBOxjHaGY0Z2i
SJ2xRuNYklOpOSuUTYt2HAgMmXigUNnVJrID3hBLlTPL93/tHfX2ho5rib0WaChbhpWezpY+nhvS
2nJ+sof7m2RH3GONUHhQStzOQqotJTcjqKBgbn8Hlmfgm3XYUqY4pjVCSlb4rh8dqvaoDVFxNxk0
ck517kVEMZsvH+aioe7B4LhiNcDcRswHq84cu7K+feanWpWFDu76KCYMzTKjK/5nG9N3pO5vtb9U
tC1J4r+QE280h0eo9GIccPH1tludVAecLv3ihKTfELuP6mgVFzRW+fdoZ32d5ruJ/ErAGy1O3bIe
Fmr8l1EitlG2g9WF4BJASQcqV+68AbShVhUOfYA+lFNVtjOjovFax8CqQzkC/nmz1Q6NWsEb7OsG
Q8Dcx6xDspRRd6teuqDcrC2iFPfpUA/YLsPgdF5FT5dI0nPibXKRDbedDY3mCuUP9PrpyVdXcn20
axN6P4Tv4voK9CHJf6J3Z3S/nrKZQgEYva64gvD4Fqbyzde97qsrhPDNOTuONFMV+wFQD3kX9fwz
zZtbo16ED910kE45RBROCN6ATLOGc5xDPjbs29yjQmFz54kJ2rDGFVBeSSxQ6IO1IfFGKBOJwId2
KuMDVs+Ans8EPWq1MS0tCGtBPOSqxiBDyCxXEdFlIxPN2FpZ+Pd6aHGsFOQuV5F45wLjtB0HKKjn
WPSNgBq+iJTldWbuKtK6UU6rdxjYJ+LD2+/mWfh55lLfb0s0EPvoTB1S+tEMF1xn1LMOMBVgwbsI
YhhZVmE5Yp1C+XQ5qSvOUySn/hp1vbnu3TubKzHdUz4eZkTUoe0PZVnh+uh4YdrTbK4tKRtrYu7b
MMw13h/vVgvathdPSeSQPrN4NJLwlEVEKU4wVJeScsIv2szYVxqxMNmCzzy7kFFviNTJJSgaH+tj
Y6OZlzpsmsBCmJY3XCaubZ61bmRwEa2kGmgzIiRqGL9caJx5+zjd9B67cMuKqj/QDD/Jon7y1Ayy
IqWw0bBjEel1vysqC4abPPOAtv4gIdUFJhfNh+SFZL8YsS+Z+B2veg1bakGSBmJtu2PhlYOYcnUM
7hzuEcUJR0gz3zWmhNAgfZq1GIYgCq/TpzscrisEkCLSdrNjjaTpKH+mmR729Ei7vYDlCtQtuJjB
3xzLx0fSs3wNLXWoOfm37oO+hgTFuEW0H5AvORG+1bxCL9Hv//oNTa+6eTx71wiwLiQt2mdr1vOI
1FqxoXGDVS0bwTSB37cRtglY6uBjYuKuZocmrhRc3S7mUwooyTqNimvYKTsX1Ga0ouy91Lu56E2+
mdeM/Ohe7tI8jsxD8Fg3iXI5c3WKHmF0rnw+OvDrb+uNNxkrQTqNiPIzlHMhoSiLy4YoLK03cQDj
y25LxFmQV6bkP7w2gbC1xKUW449SKKFOMVhtDyoOCAyz1CLWDeSIgck33odiioCZ9ZzJCEBEgz4O
y004iqxILc1t05DkRIy+UZw+G39uX4E3vlnZaXKJe92s6xGpcNYxa+Uc+ZIwgp4dyOUbr1yqPWUe
ysNPgd5LKpF0dpYyNxshE/nIYJwecd4cqbWMj33INYcmATLK4n9rsEKUHD5vVM0PDVtaqw+sHz4z
wshGs9HpRtU6QbgNai6LW+uNb+PgIEyzS0ghwI19NOYSU3TAQchB7zovOP1RZ53rrTR4xQhXvDbH
x2+1UcEweWw4mJURgsgXUqUBLvGezGTlWxrJl+upKpwbYXJBy5L8Nc5Kk5kjy2jpRTfGItsfGTcu
Mq3x4fij+5zS40ryfA4VTHeiOtBId4ppovVP6/H0c/kk0r9PV9teru9t41qKPiKzM9M+dneqvS6W
fwns3R9tjJ19q6VGbwfpCXDhPV+sLQxldk2BICb1TmrrqyARart2Ulg5XjjzTTQd4ijUtoUBqhh6
n2LNLKMBNsIQDmFd93b5CBEA9R5szD3DCbTCVzLiv4/w2fCYhb0l9/I4VKLI+TY4bC9RbRJ1lktj
5RuhHxDT5N/dQE2irb7cxPdrXICgGCmDUFmJ9qmxTlzZ7aH2MdAhnynbub0zOoBYtZmtBvmMuZDG
6q+3AsVxYV//byM7rpmfVUYAq95raiQbeqODpflBIDKDYhJYpchtWlWe0d97tHfo2l9N8JtbBDt2
8vGfaG1Dmw1gqoX9OVM8kWVOwrP3gMpmFpQdtMpLAOO16qQ14zA0CWdoXNBkvCIDpxuXECv9hJfD
CJdQit/YLxoYzt7h2FLtcvNteSU7l/qgBht+6orIHQnq7O0s5c72QmGw7tLKJAdXBKFYSQh3CPOl
JHfYNEGo+FDoqgJAHDN/oUpLy66EErxQINXtLbyrgLpa4v79sjvFUdwJ3PIUrMm00B0+VIHIPr3Q
MiFtjmjESynSAa6QurXsckNU4HibjVyqYq/mKzTzItWmgtb0DhDkQRAYKNNl8tb9XpkpF/nzFrAD
zJdec8b+esm4EeZrWRAGDH29XzZ1VNnKo6SsQzlL4/3eQU72zv3/ZFKeaoBhcoO0DhusWgrljN6W
1Y+yTKJWV3tAFkk8X35rbmF6a5TmmqqcGvbFazx+juVujtUQRkw8OeL+kHTXKTShFYjJEMXNdM66
X4EMRviE/D6XxjbN5SXME/48HmSnH+rWt/ugchj0yYbBSNpPPbs+fK0a00hcbjHq6ewJTT5GXMYD
MizpXphL0qet8dfLqa5VLbuqswG01rk2Z+kV8PXdgCRoCDchA20SQfb7O64H9RHq9rH1V9X/UgDF
zqVdHGs2/SYy+TcacBP/7RW2kH8ZncpsE/QMSepvOqDXWTGc3TaHEqLC6T9PXiOl6FfJHMdtrWhT
VSiTJ9M5HZb+vLMkVtWDeLKaMObsBiurcBCA8XreUzwOiHGfZq0vTcOc2PiEMtBv3cvscAflYeYY
55enlL0931S3ZY/Lbc7Qz8G7UjYKU+2odSknSsN6ub0PuXistpOtJlgwVmfEVVLm7boIux1pKuzT
ffeSj8Twp2m1KbqH4I4B0oi05f8xGJUO1+WibuHx5aiWTCucs85ATl3L8JoMYZ2MDT+zrHe+YURU
qno4g/0qISKNju7pD9Zddhf7Y+3pIbG9rQKwRlGVnmSsH7teCDfeEsTHprE4StoTzyN50KlUCAHF
wL9bZOHcjWl5H9uX+K1WEQM7dCU2+F5ZTvAIEd3xdafH36CGmDRWxXoJ4x2zx/0P85kC+LPRStNd
h00NtnzZ4uwW5JsY8OS00rwlW5RtWoUAFB1yQ1vEM/Pdx9/lYYnCG/jOLbuQe3VIf69+IQ2iYSCX
PunR/FEUAaybQcAGwZDlocucvtjkt5UQvUes3Blz1EPIN69k8Vyxr7Mvvn+xTOclpK2DQeRbFraz
yRKpo8LBMseHQi1hM2pR1aqXHijLlXZE6ao89UKzbxCDfpkNfyEcIwwgM90Z7AVbu4Q37N3bqRvW
0Ys8Qb6edpGFgrNvvmDSyqZ8knzxeJcnu3cnjhVf+CmKH/IbhNqWYB0ie+h+9AIf4cNHdl5CF2E3
pG7YQGzRk1eQ8LMKUqUwJX+6eF6G+mJkSsx9H8YP/c+Hjkp+p4UDhgTGRb/czgFT88Y1UCgJhU5J
eJZXbRHZVis70Nh8auWDEBm0KL9G0f7mPjzv6KuOEi/DMbu3h37uYUJ8Zluab17cg12mFD0R3O4p
EeTvWFYEYDkzO2RrLcRnJUwfiv5FGwbb+QqJAZlJe63S7f/v5cxHZ5eQtRph5EThB3wvfQvQtkxH
CCL7T0CdIkaKFxFNxL8tQj7mY9PWR75l5cB60HCnajXadxn/nWolu5s9YMPO3HEPnJ4a8V6eEklV
q5264DPQ9usCTuAkITIYFNoMjSkUQ1K7hv1PUKm70yJPa2O9KDQzE0nVZnu1H+650DIzJspMAByt
iOAKZUmeybeUUKzVrvdh2Xb+ofTCz4dBU8xJ+0OEM+kKKzCFs5NIQz2d/fVjoA9kPcR5Rfp8/yvi
nuUVl+a3dzehs5jXb/pg3kt+WnVukzYztkxncLq7rphk13dNbvdE+EayOZcobJuKjClp5OOuz22N
FVQGTdec+RTRMP8rhOEYT0fzj8/bMoUKXmBPhPJabqvv7W6b6xW4YWr7PB2n5nzlVWCGqH2S+T+Y
//tSJ8RVsJR1QpaJWek7+aj6l5JzaEDM4MIje85j9sp03VwsAg9wYL9DuPR4E2U29stZYheWfaxB
+L8KWhvgMUQmuQWssyKk7ZqDH1EhQ6jyPrCS4VSp0wPg1gITC05CRTip5gezLd82cy3uWEVFGuoA
uh/8rSRWYpXjW1ntaVZGO3JXUGZbYS6ooEDz72+XdQLtLizvEHZOO4H2+rvz8fMiKT8ecQrvABbu
Gpfnzp8VEggPOyZ1OUSocJEgG3rpXqQMCPMxJTHcfuFH+Kfpl0dCIwXaMTtM66vRmj7hf4AcfFDE
pSg2DAhmpnh6Vf2CRGpitcV8lRbDJKNjH4/b26p8xxwCTDFPDjppznbIdgB+vgY7cmf4wJEOICdk
xpXKb120Uq0TTgCeDhghvqw2fQ52gI9q281ou8POnSSEXXDeb5cpArviCTA8eOQn/c5DlwaSP6pk
PenXwjQSb/IU9K2y/y1ojIweV5LHDK4AbOBTI7yF8nS7cN1L0hq5NB8SbVQaZQBWk2q+keEkmzSj
kUziudid6MGvoxuKb+i22Z2ISoBdM9aRpuJfQP3gXIMFUJf7EZiGPZzQAMCBLIfSqA4USD3pAPlx
vDDO9tLluWL+PuwW5mrP9R2Grb8W3y9KbI7qywmvmfAQc15jdsaLOnNs0zR+kIDpupvAtcrfJizH
+Nn5PECdmlRGJj0HZWiWw1dxNoeLfFOihtPasmCillJ65QAgq5A2XJXUjeVYeKB3bcYo9G39/2XR
9G8RkDAah+4Ghm1c4gFtEpgsTkovFLVBxZTk+pTq6BIi6lMybRHeliypclQYdgb4PMM0pzze38V3
yf2AqhLU3kIHhwe2pLUyWJdQ2AoFJtFPpExLvZng2upsB8nEL7qa1AO2K4L9xPadR7xTgHxGAFAz
l77ifuPqjwyAbJsTKscKEMD3AppmPNPGFJrBasm7lmPCS8YsbXDmKESjIv50SDONM5LD49mslA4S
j4YThJE4PE8wRRuqomuJE/NLbMb3PDAl22oDSZ27wwuzwzC6LYj4KxdA74+YcW3Pwvrobd01HKDK
TGGJV/dUpj/vRM2qLMgz8ZMzQnL4AU8cgpYogBWZd4AIA/nOAPkA8Vd1Rt1+RM3Pm7NRW9UX8BIi
laPSjE4PNxRRBZu2v+yBI9qqq44rzNWAXKDhBuPrNPna3uuJJN497syjeu/dz6lFnYv/UKEv/EAo
5JjJizkcA7HQ6p+c71RA/OVjAOnd62jl+HqErvQftagAqAoFKLuHXl75GVBzjZ289vpdH93/liX8
zPVo50//6NEwT4e7Y6nYL9tQybEO2gXC2A6o+2c5sOw6mW3l1/ZjbmhZV4rHjehInNW3f/rzjRXx
l4IeEOSHpElXrHHTqVfz2oGwihrzcCi3eTj5JPX5H7EGWYnPb2TR1rlTU7g8//+Xhn1r8ugevN5o
Qv3R5ienyldhfzQUM4Up4Y5S3TZq7ptHXLD9QoCsTkc7nQi2jTjTz0Ku/BK+Gt5y0y32FXsOdGBc
TxZDCjqtUEC4KejoPsFAmwoLwUqEXLyhIVobq11vWcOSSUQh1TNdf8Lha/IVloXTAhl1NfnGPV0t
r1sSOaqpUdubvr81w2sBeQXDpeS0vgPdCrV1cAgojlMPyaWtvjFViG/xI4XXvT9lEQbOg1gz4frK
8rmrol9yEr1++Q6z3aqUSyVbE0yCqwVjpy5jD2GMuWdDEZ0e5DpsEusfdTjEnU+IY/NaTaVJeljQ
3AIXIt1h1ySK6RkA9m0JSgtZAALVhjbGMqF6bQmBb+HmSOHXA4W0gXZmmkkjL2Oo7oMT5nOpWFBA
+rzyTW9rlnZqZMsj7qa1uvXNcqlhpya1q5AJz6H8nV5YTMRBkgXiPDyAVxtDqw8n9PM7r9C7gTAr
kpOF5IOFgZeshNFEYZ4AJLWVp2WG6VdI34u43KMKr47pnBaf598TcB+mlbXM6V4Ktb+TF4oBm9VK
n0KAD1Pom6otWngaxTlE2Qh17oo6co028z0UwIeKVQ6emmTZ76PpHl3XvJjzAf8ABxrTC/8ZeNrL
l3++kD+7wo8zFDqL3pZVwofyeOMdP1x6B+TFzSSCJu2LlaKzoWCeToVssV3zoTOZWAPxGYniPpen
5t2+flKv8pbsuKmNvhzE/uCyjuHzfd0rSGRGGGQIjlXSwMoTqzthwTHV3y/HmlyEUOT5D42nyy3X
G76UyqZyrtFFs001GrHT1L6LBg5Yksf/S7yXwnkWL6K3EhAwgK4azdNgsHgjXnsKweDkHaaxJTFw
1Z4UuF3tbHb6/AjYEU63x6kYsfIZVLft3hyFVKY+M1O7JaCAGNc8V+gCGMUYO2Ge85gRj6jYdiiH
7ypwiMpmQhZxdE++bUuFML8KBImxPV0g3d3o63JMakhlZC8VtxnOMNrQCgXdtQz3AO7QnY6BqDCY
BJnp1rFNHF8nEmxoEY9oXp36JZ+ixKS7O7PJ2mwkR+eDkTa9U9pbEdATXRHdKPipGVVVER26wtD/
sOQhc5VigrUDws2PU3HPZAe5EpeRiEuSSHBcChPO/fVdFHJ+BJodcxhu/tSZooRp8zSrMOvqCmMU
uhMpGQluRJ3HQVyji9UiB+IM9Q3jYfIgCMoKu7VYqbKt1yNLtMxvcK2nJYXeF8ZqUD10ObWnugHb
BMLHCYGHE5/kXGfqp5Nxyc0Da14s+apfTQGnJlTTz8dNfgkYlxYL4mu50H+j1Lz1pnI31a8JgI2q
gaZtPmcTh8H3uM22mEWwl4W5YALhFdWhnHAW4s8ROvgOm6r7pmlN0f6oLquplliMN4fFycgq+JPx
TIsSpGaGq91TeKlX8KeNawvznzH4ECRw9F9KXcA1x65NhSBY+KEHmn6aIrtIhMg15h1qozLKV9w5
PCRNx3eK/+B4yMXA05TneEBSufoj1aLqg4LMluHiNOLJKGU+CO2SoO5ExzvscwfuTxH+9UxPHwZ3
E1Hjnga4fWXVudRYkHsU8bXAFlIG5+FvVXOleQmAalfnv27Xps/O+TcxaEmcbIz9fKHgUFnaBlMg
Nnqc+AaQmbKI2GW+HRrKZURVEYWdh8pUPVI9W8EzFyfjl/f+KgjKmi+gGyFBQ3Dixf6cWkahTrGl
UPWWe12taHwiUAoR+hm/hZEXgwKbvDg0Cmo5KtBK8y04L8kC63iMPbc9b7Qd10IKQxq0aoe5Y7h7
atZYFIff6F9FiWWytjT+WFdphl4dquNhpdyczmcPa0zLqHHw4afiQAhPIUqyHl+2YxhM8GzXVMaY
OLzwGGt4Pba+lYQg0ksjFw6Rjv00CGVS0b9GnVU6kmcvayg0ZxE4jiOl4hEWgAVAhsKiFNDp6TxB
cflX2mlTLd2cK4G8o0/SQ8WfnOBB69RoUu4wD/qdmd2kaWZXdKDxmfzrB+Yye2j/jBFIwBl8wOAP
M08VsCSoM/+nt08pguc150/T9sfCyE7k+8GgyrfICs5Vet8I0I6yCLDG+0bal7yRQLvapORKHVwC
vr6ObtivEm6EC0SzTFXrhkr9SXRyCHSY8KiRa9QQTTbg7qeOBUVFFzOtpPbpYTnBL1oRrGTa1yTo
u6ZZ347RdclvfsVtkY+BVBouwooJv3O/Vs2zEwu3nZwI1f0X4oTPDuUNfJj3HWTjY4wsAYBUigIq
RrbdSgTI1AIKCWspV95Tc6+YG4DIkxh7YLt1nFH42ZJY+35vP7jqmtx6pcgYVG/Tm7VBToSh+a34
jEWNnEvW4bmFq2F+cdvoSzPWpaNtv7oEuOKzdGbmI/iQps7ospcY0VgMQamn4CkoI8EG/Ce5Xcrp
69oxEBUzCUHzYFpZSRlFYohU9udfsGc1rfWXYvBrFwwT2ZRBVS7nkt6RVlVl1yJUymuBWZbBpTjL
xOma4fn7k+qfaCxnjnpOxO7YNt0BP+wHM9l1u9gZnFQgJfJyYnMXyii0P97a1jIA8+8PHwQ6ecA5
lADpHnh7y1OG8YyEfXWM4VNrxopdu7/aL9TpIA1dHi2UrLinLsQ8zQeUhX56HWJEjNBBZi55hVW3
WkxN1aWKGvGD7oXhpB+VFlZ4GXGodBd357A8WYCKO3HXuAlNV/MPV6GxFQz+ldbn2kvOKUJ/Jj1z
AJnuOK1IlbmrtmQSUePOBtAdV1yNVLmva3TQylLb6g0vG1VnRIqSf7t92QS/s7/WBXY3EDGu9TJO
IXH5OCIRhAJv1imjfyHQRJINS7GG6vq7mZLfLuS5sdOrp4HbnyVKhUKi8NMa2j6+qAsxCjfrMjB0
z1Z1+l+q0ig5OtIDZioSnTIqAJz9vW3fd7B54eG5muIOM9TyLWtnHXpHVzNNFhSKR31LN38GU1kS
l1wsWdYBOXxI01TAurDoJeXHNt1Y+E3oQxQrGnhq9uHh8vLKBxkRkVvccIiVahWEI/0T1KsQ9JLi
YrSZpS+Z5RrjTCUT1LgrBkXdTfHGlZLxAliFiQ3hKFcYpgzU7pD9bMLfeK8BbUvpS0PzSbqQjI6p
E0ziDFh/BW4Pe6RZowQrLgi71q2gmDRrT9EQVSJ6Z72ve9qcsT4TMpsJEz9pxMaoPq7Gjj+WvyNS
/z3dCLtRLZip178hVU0aMjVGwwAfRnJpHhCo7BxH15R2JR71M3q/CdlIFjoQXwgyoTyviyGMWIMt
hAb1uPkTD4VFWDAXVmwFmg5+vgh+2S7I7t+WpILfmdi4HN0kFgzocDnaeVZWbG2A5P7jIaEX9oBk
bk9vusrZRzVcg60AmdCEin330dHcMw95C3Pj0zUi+v1Q6nfvz2O1RjsshDJmljCejzqbssvZAnbF
WwqKaUHwfxBQo9aQiDCEVupgaoTuB8Xznut98MD/IwjeBKnf1CHvZtau3ybYaK4qNCVt48ZKr+co
AjTHM1Llh5lblXix24ZDbdArxlM/YEU3HBG7ZAhXlayQCpef/E9fHhdXxE9o3YYgXadP44ZVwF2G
q2tQYi/Ltg2ugJOe26al+mFlKv6lP80ZPb0G6YfS5gHuXX8SXALCBOiLiRuvIKieGfBzOyx9uOh9
mz4qa9IUGABjqwKD6hA7wfkbmJioyboUFoNZEaKASXYoj4HDJzBRMlHFkNS+DCa0RwkVeXC7HQo3
mfAce6p38DRSpcOYjndezs7K6e4x2YHfWHKcgMXAhc2lHOW6PRcEMffC6WqT6o6o+nRICCAZMsu4
XO9Q6DD9XQoas+T2gUo7Aew8oGyqdDFn0hQDtIeOuP8N9bCbT6JEm3GV9lMpC3xWha0HI3bMNj6n
zF6zqTmiwPYOfhWdlp6MuBGpfopMoh40sAIazT9pDwWAQyV1DL+QqcWyy33B8lQIc3RHm/cz5p8H
U3Cku7feQgJ9UNEh3rRocJOcGpRvUlfFfkd9cyiSrzsOd6ocnck7bQIB90xuiAA9cHnS6rjflKxY
W0h5Zp8CFq6AusnRGcjPAPI6Zirih3HE0MImcIirWRK5W07M/fQi0oSfzyjqSiFdTyJgglX6glzM
MsgEffyMYUpFmmdUDQQlxBIoInBAsMdyfv81Omv1oyh6aZJHHPfooDMJgg2EySBWz7yTqEblR+Cm
ysksakdpzi2RaW3KrJPZJmN++dwmw+IKtbWSXLiR4oM7pRFmwC9swygu7qYKBMjkl76ZyhTV75PB
mEZPy32A9XTV0DpnjZcz2ZhMCVmeb6utc7iQOaVLML6nJTP1CyfeZCKzb9r+OhmxHOwZth9nb6wI
YNTeaRHBVgMguysnAg4cTYeAF/UACsNg8zqNps/FmEGIIPe8wmaFXqhsVjPJzKZ7ubur1v775Rcu
568pOFb2G8gH9u6WRTt1NwI4WiUCZzCn0nJRFEUbrfiuP15x7LC9Rck/IV8mLmt74ysyn2IYXUt1
lOgwKjUuqzSyVmyR8zDWMiZ7r6oPRDYwHqeZm4QoxRNs4GBDh+eQ9NoQnPs2JjrNTeB9QkdLTl/3
payhPuWcuDFX5C6N+kRa7PEUiJRPamMYpL9NwJzx0iO5+OYj4lrxza5eeJY2eDxCVCtqgVnpm4or
4K6Pr951AE7yM2oKKMV2mB1phyiO2TCcW+j9AxlJxkWd4zahm0CM8OgOYCebZw3Prp94FG9cWWal
i7rhlueFMECPgLU4PP3NVdDcPqrZJfowCnDQdOGgkIcSe/+jGQOIT7ELRXhUC7UMXRGF+JBk5nF8
vqjm9d3TY4hXEZ2tXJVAp8YocVvff00SLDoXFx3iv5hcby5QHhC9DK+LngTfm6AHtrWFWzXmQlc7
SLL5gUYeaOaCOFVEhLrU9EaGzuB5xfrKk9fcGIZ+9SHoK1clmhowJFTKsq89+sPJr9TAV+IcxM9+
/ZTu4TQ2aK+I2SiT7jSzXUcewwl+fD2svXW7Pi3z1/g3ECosIq95wRAD04PJdeDbLKFn4JA01OWQ
eq3VNa3TolyCrdQ7UsWN6zw4Jo4Ce7QJ9Z8jK9bb32p3nl0EipUwdIwgmTvR4UK0eZ0xR3J/SCVx
9hBb8ua6UZxTT6dgxjTBVFAbJuIlE2HM1Ge8MEKx9H6QPrkLgRtFzCT1GlyRdPVKar2WuV+KYIXw
Ki06QPm4GcnirLCuNW9hMOLJzV4NZwc5RyAHsRAAde32hVWuEcG8cDrr/Q51iTOWXLf4vJvRQ9mW
ZVIbWgT5sElAaFZyUNHQHsJ+FzyiLcWQKN7DLStf+bpsozAbr1PYWivRhKM1fTAlstQZqeaL8Ftk
ZKWcF/EgLssB/iXDBztBbkBfKQEOHdiJT1MgZd+EJ+1pKnLYhryDPEBZAseHETLfiQ97Q2+Af+sm
J+JBTK/iZdnGdT0niiRzG+U1eocKbZYoAFxdBaJjryb2H8BafbNt0sXFcXz6/vhq3OGz/HVyhN92
AwHbppDXaw5MsUYPhgKe8ijOn1I8U3YU4jBtM5uESCOIoms8A51vNT3G7pUvg8q9LGrEQjEP0BnQ
b1tS91yoNe52yu+B2KYvDgiKSWNs+eyzDL8PYnLWiIllNvlGCuEsI6K+CVxwl3F9UXtCad+Jx8R7
2BmUrpx6f+doCLfnsRwiAJ89VFmB5U0YZbo8lAECEqvOw00q8wF92v7tHX5pGg4017eeGISdtPA2
uq5TV7xNIPTAXyNyocA9RXyrsZrT3FYQFyPl1AxIS++fi4Ij3yoZ/tz/ha732VdklsQLalS8Ue5o
dbuwAmV2scUAewtr2lMn8gCPN3FXr3IG836KxElBAqxfmSnF1IIkaSaotI5x+Ob14XCSFweDYXa4
Apmecvla+sJNKfNQid64zhFFTFD4cJOYtd8Q8haJdf4Je/xxqkPEtViz/PYzQFQeLyCrP9GHdYOy
EwBhlzhlSGJoPAXtgYP34YqlX9O4jUiXJkMKtTLflXXGJk2FtTcJH0jlsG7kUXiJWYaRsPzXri4z
LzfugLdijj20b1JsDteqedYy5thggIprWOKLji8H8XfeMjuGItTjx4V+n2FYpxW06T/X8l1m+Wvr
QdR9Iwo/i6tgSUQDaSwlCBW6/btL9HGOzXpI8cxGvIhj3iqwxNjJ1Pm6EhXcmgXDVGILzRXJ4NRl
+uOmXs+81Ur83ojYrxlaYbhNC4uB7lO+i3xEJNe6CwnoZgHBX9qMsAyohpiGPg5bivzMgRVWS/iz
2e1kZkJu5h5oP0Uf4df/73s8YfgU3+Cl5YkIkW9+opxyJITBygLXpP1SOqBTfivLK8NMuA3RW8aj
HBRrHGlph63Fei3z1VqHkfUgSh035rW4E/UsiFXAmdkF2359vmxk8EomtBR4NwebY35+zB6LaqFt
9bdpnl/IdR846s9BBdqSiAOFBxE+GkZGshWnkHRfhQKM0vrWmHl55BQm/8mULLxM49tbqbzF7Tfp
uJfikyc0HAcCTOef38ScVcX1Zu19me4aJ+AJli5FfMQbx9Ifn5WJnY+iD9RAuAidOU+LPOzwPg6N
uUzsu3DGxsltqVldXDM8G38Q0bA+GeqR+xIUlJz11NueEY84JTPEVyQDknIvKa3r4ZJasDlg7F3d
aYyLnhVZ5vMGXJvFDVNCaSBi7fYizLUxxgyBc2BhLki8l8Wi7sdubLFfKO+o4+s6Uq0NkW3DcA/+
gU5Y460e+3zl4Yt7q691Hrb/Tu1/dtgZVLNg+2eXpXK7GTSRDE77WNTrcS3D0ovhqmCSmpzgqUSS
efVzPa5YWlKr3DKvEMj+kVW4E4BkFA2U17hDrabq5uW0EakFPUhzLxLweNLMI0gyP5LS3dnQydfh
Y4Pyr0Opx05tT/QPgjBEdfRIDMkP9mnMtk99cTrWSi0K5tutZSSZK8sSbwZ4DWRQZmGdWqY+9+Rg
SRO/mC098jp31uMy34oJ2XNJy0lJZlD20XPUPpZv3dtLYEOFXtMZMBL8nrZUHrSHYWBUvkcL37Ie
Ih3YahJg9sU19grVIKYmhcXChstdo+Tp0kIUkRtxyJ0Dqnh/pKy7ZxMv8lvgi0BzUagZY13rchGL
nWr6k/dgjwPoD0CBiQnlblKXc7kNjQuSSeoR99J+zec2ubbToYVx7dBsj/KYtrTSIvz8azLNvf0I
cIYu8VMkxBkvXjh/SDzLq1WwG6I9Whr+wePf3SsJKYlDbteu0BR+91xSiv6hPR88aM3daF5dzsYX
qTMWdQRFFHqj6IS9CX4htwgdE/1/SqYq2UtOlSPxc20d/A4I6ZPAbX4RY4pEZGKsFEsyvaM5IVP6
nEWw2HphxvzzTcone4JFhdLYygPcIVf8C9L+TflzsptZsgKvl06XV5MAt+GoZhU+YMS4BPmQnHtF
y2e2Q1sriVJ/+q5W/ydpbvvpBQ5eNV4yuIa+E4St1oqq7bY1yjy1qNjXm7IaJAbL/Fg7y+9Ablx5
SZWyyZxxYuJ8RGYPBRw0zzedQu2KRJjr1v0JrlGUeX0g+NvElO6mxwfi5gFvJpycLkYJUYVls1k3
ZawbrH1K4Xm4C/kLB+itFtRkdDzY/EPT14ILmnH9RJXu9+i40t+k9G44SVuwMYh/jriP4jbZPfIe
Ac7PbNwOaeAgq2vbH1m8+RSKOyT5s7NmoneY561NKRcCLSajHoAamxTrjMqGO4JyxMJar2TGhxYO
Gm95+uQxRp8J4OGaplOaSVBKIfKaRPhPDszQ4MCmx6nMjm2HNOPslVhRK/vOoGEz8CzZ1gT7N0No
I43Ar+JQAAeoeH8BeHRySHzE74T/Tgd5WeMF1cGioyB2+EYL7gMVwn5gfsenYRkAqsd5YIOR6AOk
wfsNU0hJnvuAAoXNGrQzosri7e4b9tfeX35IENnDNbzyNtvUqjDFB2+YqmHOIk7c91IjD8yZl90x
5WA8/ae0n4+FuNxxtr4CKiO9FE3LOc2aNGFhfm7irpiWu+tamZmImy7OgKwWuN4w4fmBjdgpKpWD
/ZQHLdJlL/1CHPt+cmX1za4mJOLC1OtKiDhtzbW7zXzccrPJMlaGnq+oFfPL7xqbyiDxPlQSriAx
sCQvCNMd71RaCShi1vds3tNYu7qgUuNiFClrxkWJhL0HVeB/d77X1tGZsaokkMyXinQ1+hLavJ9t
lTNFhAPJhwHbw7E+OiYhhp8pxYFxpSJP6g7tDYFoD9t32dZR1QM2a6rzgvKSgO14OWbAtga7/pmI
VbU7TeP+aLxf80daQu8WGPeCCtbm5A8TEgLSuNRGFRkIN8d6jyJuvxAjHIPgjUCqEm8+MqsXTNUd
98kjOyWlTWTMP23qJ/AMaW5ZCEP6XRoe2uYBH9XobTguX5kCr3OCm1Awn/SJ8tXOvNxCChn5Bf2D
fO7h9i0TOQ5nn0KTxt71tzRBav85JoPgAxWCUsFLRCG/9V4mVmYKHSkgACgWovsoSEY5VCkLp3IW
4xUnQqSkEI9vxeCSWa1U5KkJm1sDUBC6878ZSjxFDo7NtVugRMnTiYPu+x3Dz07ujzWAAotp/R5E
2SNlBgBe/vK8hPbBxVwDQ10DlCxwqHxIwTnWOgRO5pWgIyIdpJfb1zcBVQPnhHo0msI4ChkONJ36
dph/ZF1cV79pjYVlT7ELoYoypLV84L8VjFaBGMQOeBDJv9snYRyFfWjaJiSGeDxwhhJsYAvCgRo9
5+PnwGN5Kol+jAWPEi0as93GerEYNBmlHTqtayo3kDURwF72tY2WmNUdi2kl3NBFbAsnMi5nemis
aghA7bNf+L9z9AL8ZPqSQLP4co9DhXvNRfOHgK4wQDBF5Rwn1sDwRXiVGLKLzQEn2MzV5WFG2+gQ
EEy3/yioRqxzK71c9yPtuv/lu2vqm5DyBpB+QUTQxHnkq+sZOJdmqqE3eQeRiPRqZAyq70cmDUXi
QIMlpbEH9/QiAAe3XO5peGJEDx8iek3mx3D80IeJHHnl/L6/lhVZ+ukoCTV29EaFCrD2vUBGmiZU
BCfJvwHuSOjTMzZzlgedFpWq9j+lTMhsmVvwXnFbE73ybBg7h9/yJZLfaQTAWQWkvJcOhYiruaYb
UZIBc+cMFV20gfcJhalFhNXOBHdHYPeJyyUjMrwEEVIu3Pe6an95G0YEEiNepi85tAM7vElrEFRP
3iueWi+edECPYE1S0/bABZWVJNn2CNSfp/rDXiqVjy18iDaeuCS62kBgfZ2c044FPOb5ZIMEi7kf
T76ytGwt/AjW59pobVnyp8TvIplyTWf82DyqqfBy0weq6h5HIozJA0aLLHSDlN/mkV4MfdWBbeyl
7ii31B34Xk+kHMv6M1z1iOnL7lfVcMIBaS03Hijc77wDNFkxAa4Js4KAE6qsOPlCl8eJELe+BVTo
hEKXIrRBnCeISkCpwx5eBRCQw264Fl0sMX6OX6cp6KRRUL28osG28kXagmn6x1raseBAIpU4PtgZ
u5ldMawZVW9qqkPn5H13Ukkp7dm8MImtm1bL+Xfz5UA03tghlh6XJyYCOuLgy9BX+hSd2aITXhsq
j6fp0+/hIuePme1mG+EDFdUijbHmnVkb3Acia/7atC32iVjeOsAfgEEjf0kGdvn3lmsRmj5JZcMG
7uyi662NIqadFtI76ITT1c3glUNYTmCMLWXiqgA6S5IB9EGEKra6aWv3V4QSY60xR7BY2dc1Ivps
x1wZdAGWyW1x2wLy9Es/Ns0POH99owS1b1HUs+HuSYRfKsnmr1Rj6ITY9sjuejfdeP4/AkkCcp8x
BPovFrJ8gzNINwit8J7LEpz8+1Nx+ueHpBIftv/B0Mf23Rsvq8NPTK59RIfjNGjRDFgNUOJxnc2c
tx/GjExqTuAnrHhmS5Qynwx7offaWx7xZrsyj9TriD5Jh4BtNivuK511eEfcvvwC6GGll43nrqB1
1WHiYe/NUiALwTKIwGKXzDVlt+30Mao0K3tXmziZLaa7YM57DCGnUsgUkI7cNMVpLwtTNnK1GXQ/
WALNyUlGNO27av7ItTtSzvivSK0bR7AVIbk/CfkQLeceryjQcQqhqOSbeLvqP/RFpX9R6MT2cA0L
NR5CJiUetbyiAo4wOrLKbls7luk/kiT3BRF+l6eCoLW5Js5ShZtl9NZxNCc6Kc7jRhE/drl8VPjD
opU1BynXBlMqT/wcRytPdtE5LNzpeji/Y24LUqBzl6ZdTxYYf2U50p99HKaMUlc3lXRMTD5bXzYK
AHxkJ5IjoGCg3VmL0jZcGApf0o/n3Aoq39sQ/3DbRxoHk2T+hugiRFR01qKvzX0Woc1XXxVZx+5W
ywtbilwhMtLDVmj1eJvZd3KzLGczB2lnQWz0bmQlAzm3whKtkVK22QJpSUAz42aYxHWSpHFgQI1H
cYQXjm1GISWS8ssjuF+3QbFrrguNbyft16W+xfhsIgx9Vhq2CgTglmrxcTfA4T6dzGpsiU6y5cLj
6Bab1fixB9GykhZsMiZv/AOnXnYMLNiMP7SSvndZAe2GXcchunVH6RL2pXpACnUY67jVBYWZw8E5
DK9FCCJTTr1LcrarrXOqp4GwIgJ6qM4xaAVYAyjT8Tusk6EtfZp9CTd8tXRKuMemL7iG468JGXSO
q2ZR9yX5gnu30Nzn0adn4QOnpmjMhzotr605sPhG9jkn+wrcy1xJ8mZ+x0Mwsf+/sIJPl2lAyGD1
FrSwEnFQrKqjTGX6tWynzIuiJG+XtXUAlc+sZbnjtHwG//wJo44fvZXgewJbLsnPMW5/A8oZn+KX
wDQmffN9NZcZcPX58piXWKvxVMKiS3V6lfRiaKv3mP7m4SxPl2Fzsgf0Yr9mBEs0S+Bfu5nzQTOX
6ppLdjeZ/TQ3b8Ma5gudrfREVX5Tk4TBAkD/NGsQkyFBGfweoP/Xym176DUFf7rcHwhBLaafGWQa
jwwj7s60R6pLC+4rOnwStApOFqLxvEMw8raBt3rOO8pwWM3DUMVUV3DxUcR4L20vjsvn0HVEES2N
NYmCyfiIr5roSyeb8yg1qoGJG5AuW4WpzKD5O09hiAQHOm+9Rx7JUdVWCVCSOgdjbqU0ekltav/Q
ZnUEUGCkWcLxUy4c03WRogipTCt1LISU23T2dMuToYZbpMWTDQmpREg2KnHWmpWKAxeP4ckkX1RX
ZdVfBjhLMf0OXOfPZnspweupll9O5IbBnweJbkpe305Rs2WdZtEw+74x4+81JQ4T4lcbqXjb7/SY
ihGWVBjh32mMT/vpGkb4RTbCtueskh0TeJJr5jVjJMFXGqI/bnWVQXOGdPkIsIAW+Hjb4sozhqTy
I9+oY3JcStODqpsl2U6JIBXN8TKSxvi/JcIGjqQdnnPP9ifAj3eyxi2Ap4o7Bt+3R5x8O/6P9OPC
IB59H9Bl1DwKUoSRXfJGu1H1a+zFGonZNiDIG1PI0rxtQa6uNMJ3koEj3t+QlSpLA+Fnsfcshv0F
G7fCIsE+v1DjhWDC4bILWvHvNL96yMZxgGA+LsiJwBCRXctT5IbSyJVZ+tw7xXjgF5B18G32PqfZ
RH7oXQ+nPbPK8Gl5PcLeLdaG+Zgtatw5lVOUMyaDWVt3zHYBM8xFTmFwLk4TM7gpdvx4xP1H/yoT
ddUAMfeE41A7IOvfHcuqCjFRLyYFF6zOvhEPJnfCPbwCVN4RRs2yyzaylyxOwpWYKW2TtY97FST+
xojAtrntiEy/xGwjddEenYBTOSc/KjkJazdd2n0J0fUIiDDbL/yPaB09mNYSGA6fVofsLFCwMJDD
3pqaXRnfN8uDmVSRAVYF3QmsXxfU1j6iLjO04otfYyKDZskuYZwafOwAXiydK/4HZKMrF8kv8qNu
XjZjC14jtTxbFFkQsAUMGtOaQaBsy6gHGSwQV+jk/aiwvq9OJz0gkxc7awi6p7YvcJg9BawgdXxX
5fjKfd9VciRzvWlQY2ejzCzWT/+02TLAjYLK1BUp0IWiedZi5EJxhCihjRYFyWd0Io40qMUgtDqU
WgEcjhTw9fTKYYkBQP0uWQsmgZibHj5CVBLLon8F3KWBysTtb+XkEZNcRms+s5RnCp42Mo2xQ96B
PE+TV33jO4/PJn9GUwFUDqnXxeHbTMC4zfaK1gUDnndj7qQlF9/jWBCmhrv/LwJWR8jz3JFNNJ88
vWc58BAyXyGaTk98WEO35CnygnDTOMUl6ajNb598qoxChwudIW/jteCf732k4c6qbItOnYreG/Vn
1xdoipRp2G5zevh36daHbVwbAPNBgscvwA5c/AVFKzxG1yvgUjxbO0HmXxa55aOVIL5gTE8ACCFe
Elf4LOIJD4y3tNcMegf3nwKhZPp6wOVBDrP7SlXMf/bwYa08SdIVZlUcfjXi1XKaxZhGIHmBIrvl
TUExSWFnwS31bQX0zurXWtjcVaf2fljPnebmoIFIRXfx4OpZS7RQgMlm6RpfnCAvKkuR2ETsMfmH
emSlgAFWsxskTPLSq8sPKcCOw77Qw5L7ZtY6bMryBHxZ59t5xtMVr6WNtZDaBr14URlqDmIhu0Gl
7B093L2m5798vJnevHmubC/fub7cOWuyPXnhhTVwYmwCSQ12fg6fCHrWmyyCG6QZB6HXxJUedl3s
WAFfD6UgaaRqe0Vu+AqG3eYMR3pPNPkGbbYyUV1BWLrYNZMXe6/l8PEcLjIz495w54z73DGOtiMW
Y1U6lA+QMxSmOGWDb6P3ni8+q1+QnBkWdI+f4kCvWTG32aBhphO/cv1RRWQKVzWnCF2xRMqBqeN4
N6xuZ2XQjea+tieybmVHyVlLnMIrIvtYA+zNsDawmhnyomgPFuMH46VSOPbrtY0Q9YW5i6B/4/vI
RHrkF3GwdmfJzcs9m7BzYFyHTJlHAqjdWJswxx7NJs9kVBETaphF4czh2uHbRbdl720mzdkv1X/q
wnegHFf/XMqIrOAtpzc/eedpMdwNQxZGi2Bot4/oKw1FDC45/yUbcg9NtNTqUYJxiqDwO9pLVjEL
qc4iGXdvp7QkgsbtMAWmmTE1gUw3h81w/qU0knG5Mk8S+YRrbD0H3PAwxxwSWN+Ehohc4G6LdBsM
dDu5l/94BxFSAQssfO9zCT5KpPhRWSwpgjZ+8y0CSt8bgJIAawhB6QrsEL1ssjxv+ocAvBEdj6by
pIigc+FMkw9K7MoNHOCe55Q/75HqEV4nMDveYUwOF0fB0uGYICjZuj6rw4J0BqMHj1gphqK/p8cO
m7lXekmZE2YgX/yalomvDmmkXLgb0deDa7iv4aWayk72Ac9psmUdiBKg5vNwNxwcxyscFBqIozcv
s/r2mbUKdMbNrfh32i+M5K5Z5awsdh5kayuINrIywHdjSCnVIbbfjr8T5bzNoYjfDGl22wOGHhfd
gSDqkCFMnfjGb7FH980nnS88hBqYEJjwSZN0DrytnS5ocxQVBaDLlC0wlzx6rKHtCd5qCvvAqN/d
5nA0qVzzsqd54IBZGoxA+g1z9GkXrX5Bf/b2qVxe8Xtk7iwBxotu8l52ruT35gstTgx/R29E8Lwa
jNPGp9bMyzOybDROkafbXuNd4e8WZ1gfJZJaGt7WCKFtP9+KtxXUyeXALhoTrARDSND7Dhv5L+2Z
uT3ISJRQ80whw+YJ8jBWnIzDYTnOGQVLlwFCik0C2bikDxMqz2pnvkCa/Ipc04t2fXLw6cbC2PCH
zUcTGegdbO3QS5RBFWCrvMA2auEbrWXBkJN5DLB9jNWusfPcCq88gl/5BDt1KpQrCHvwBOx7XfY8
gcQc3XxwzWn2Wk9zL8cYKhM1NzWfRHrIlIl8Id8GdU9VYD4gn52mPgnwcNjmom+XqgnQ8HRyhkt6
pjDl+78K208CeDFkzibYNG7S/+KpZ9w3P+6UzqR+V9IyFYYUdX+Pb6sYUwUtDDSIVDvydWucJP1L
BPf1vsNw3dyjYm3UGHWJA1qLOgbLNaQAGDeQx7qYkXdArTMJY1pRs6NT9ddzop3AgCBoRX5yLWoQ
Vo3DRsABlgPaKyebjszG9Z0PcMR9Wg5P/+nB00HT4vGcwOYgnIfyQKMkZypnOfdjfsc49NCd2i5N
dMcATvUwxLY/fzt+urX9k3EA4iFa4K9aWNzNaczWybwVHtZsa0aHf1ZvMtqaoUjOeEeZG6aYP+/A
5b+6eHAIcdE33k8isFDY1tLfccNq6xcz2RSTtwf06vyU44LRj2uGcg9lwt9QHmJpoPSk2xoGXEQb
DUQdDBA73ve8QlFgtzS1r/f1yqtcciA56jIUBNahSvzIY9odxgXjw/YbGwwOd272FCAFeXNhqS/w
4orZp8xYFBfR4bTynn8WGD/2FxVcLzG/gsX8ktVoun3Ami4p3yS65Vb9ciMuXxQgfnt+WQuYL3ws
bhptmHu+Km6ZHRM1wYpp5fs22YsxIjxlJC2eVwfTzb46Y1vy+1263DbuN+1sDYSq3JWnf5QFowe7
D2wy05ikwmHZ18aa7Ahc658Z2mkpsWpC3NgqEC6ch/2opHAgOmm3P3vdaNXs9pjpji6veR1UtKZ4
MmM9CpczWBKynf3sT+RqxpIaxfvgmXFlCwrsSLuufAnSTEoTEQ+wlkkf1Si3b88BTLA2GVC6NO+W
XKZntAwCBByQPBbywajzW2FPv/w7/6CdK5hH5LA6V5jELEt3UQDZgwLHIzZaEvei+eM04alXAwsw
IMG53BBcxKuyLjYqFvhy7uEBBNYZibNDVj3aEGGrorqj1QCdz9hn3HDw7iSHsdDSqPuUEVIx0NJF
DJJMnmt+TXsqePvmLbP84bPga0gCuJpCoGorfuv+KQRnfyHDQqv1qxEcS7/TqoGJqUPLnCZPmmgZ
ZnUm0dERtMxHwYC/M/Loy8Sta0qX87izBrIy1gC5iZUCXJ5yBSrY7KCsbSlzeoYeGo63lOUCv29b
6mPaeKOxrpCQWK1PgwfSVUO5at99R4VO/eckYLnH3lqyIf1vSu97uMJ4hKf0tNvpXgkupGhrQcUP
dsRQb5NbHlFWg3g49sifUy9lVzhdHJn/dUU4CIF4iQDIJCRQ7jqbE++BazGzK2CkfbJCH7/Jcl/Q
ekNKAfPMp6THItn0qEOhxuGLc8tRiucV9GixxOF4YQ7uGfCdtUIe7OIxMmvJy8Qes+6tUhP75xTC
t3NKRRmLKAT9u13LYr2qXjQyw9Y15dzO3fJz7bJ3hNdsXJaKZvjEmvSsXfwgmO3psaVT14G1n68w
Edd/3mSZT60b0YHYu0JVHbwVx6Gz0VawHsTUMBn6r3mQtYxSOMHGlgPRBBPp/4sqgjWAMhoeV0B7
XP2Y1lccJTEyKEDTCI7CUz6zT87Az/mZ+gx8A7XfGDZ5bWSRJp44z/HRR5bwsfWBGiWDyDH5LCLP
QR+j9EQFm9mVZzds+wCmz9kWa3G2Pk+qFwWSATtV6FV99IvMGw9kMJby+tlqHTl9mgedWPwemXke
7TJcgnA/UorNRuFeGK6FhX+cpJyhGSscqewt0BayXxF1/+g4GxPeTInekLYzpnKZHeh9V38IlxGd
sSdlWWzmipttv0L94LQFvDAwLlezVhHQfzSZqBAEuAZROBaIv21VduB4EafYQSVqLecd/DxcbM3i
Uv5z9gvyoLwa6AQHuqOp01ozGiKTmGEn+YKxaXaTfsc6Hx2mlyR4zm32+kNGy4kW6WFgHpOZnUtQ
lv/HUC1nSbIDzj0LdVIjpIXPYdexNqw2qoax0SFVBUHm9vwNGOtXYt6wzYeFbVtYvQXbjLBAzlLC
Awcr5vp6qqvkY7ATOYDr24WHZ8WYo1lCKjZOnL/k3uvGlYDA1VfpgfZpUkBPgNQCydTMBJVDmqm2
5+xRHpXVs85+fzh0NF7pWdQUTrdylAhYdBJ2Rcz82746D7wam3EFFdpRw9Q/1UW8qrfVEa5MA6LR
rGg6gVay1oKVv1dNl/WWp9F2a4NjQR8f5Tcao5IO6c6k3BQpV4ufRcUf7iaiZKUgwFlkQ3w4lTKF
WhchtN/VmjEodAJlTh9LX8eKORBHWQbbkecKnNj/F828SbtNqnz4q9JuOzyun9KhizV9E09Wz9NV
jSlNg+SP3TGawErOUg6BkHGt4ZWsj1opCv176CxtEApygCQiVZGF83WGQpPP8ukM+0LZjN3+oNK5
VD9KCvu0eiIHk++w8Jdji6We7EdSf+PFai0B6VLFPydCQuQPkUSvMl/Df7b+HGeHqxB/6ZgRUcN2
lHfRzW5HwCrUKPdqpL4XEaoImpvuIVYCv9IN19KKS1Psj0wVpxF3tWFaHdC3KFCx0xcNPbUm3nul
U9WsuAuuJIYJ58/QqOMpeWH6uGWgZqAxiVv1D58ZpxTja0YiU2OJOsfoyWb5lIEtfpdCWGYZwO4/
DkXhIyIuqrKWX9jWlh2fWDoFauGPUyFIfsI8OLIt4zUTUvMvQcxbHmHt5QqdrAUKslJxU4xIoWaI
ZTWNuBuY82Fre1mkucO28PynJSSOjajRBn3jyaaWizUyuDUgfVMnv8A40eYU/ghddiF3m+31j6XX
jfJVQXda+ujcIiN/2CIi2GtAdhVHZUbUYHFwME957cj+7vOeoYsC9BRUVG92F2U3dL9SpGrOVj+f
Mm/naOt5JPleF84EXLZQ2e67yubNxYGCpQHwWpW+ms0BLCNfsDAVa8iLQwCrpRQhpqFIPB7uMKS4
kdYwgi3IFZ8Q0h1lZM84NDKdxQzjxFOd0t7ufqbyLEAjZKqxOlx0tYt8zjjv78nt/pWMqBZlMkEq
IEW6QCq3AaeXvauQ5KfpQw7Wg0cNjUEGrPN2fX4LwUInsZoZoiRarCthF34c1kQkLS8AjeiQIWHc
JL3si6y+J/CQC63mGjtAQytobF7T+koqPjy9UclpAmdVlg7yu2TlVEZKaUNe5TRL6XomJVMAJuBZ
8DrS8/FqHzTbrpdJlpfsX4Nemok9G7SlAuX5j7wEYcX/mLduf8zUAQp3CkKmjsBzvsLa8meMs4nJ
k7prYf19AqKXzCI8nOTNo/bZgjVpXVPQOgdlGBHZ901Z7u7WgdDzM2MNgX8rK5nHioXKHQfVuewm
Qp5oKrl0G7QtTas5VyVqIdizOpnZxVizs89agOuYDblpYfzHa/ZeI/vWA3rJJPna1lHd/GSr2t1x
MnW9T9jTUWbbBL2MfRXoAHiJvr2bJtj/IMASKvECB6V4Ojaqp81RSj4N6snkG1yLLHvh6l3GuM6/
tUa2x8SwYvgn7jnrqFDApbT8QvqMsDlGkgu5y4W8RgglOIoS8GfqaKv58ok8oZs5KV/YN5a5k7zY
DRVpWFCqnscmZHTiANJXbuOaCxK3EslCQRd4YDa6Z61aYICk3IhL+lRrHE40dHmKe/tUi0PDxi+O
UjJHGqDFe3Pt+gaDOcmr5A+1zpWgIrf69B/w3uOwNa+sVAtsjXpFlkCxhmxyLlgFRT9x4ZtO3zp7
+MTSAMYwXm7otp7PqCgTqyziapMHNQa6asxCVUrOJzlCYzAWTRstup4nDfi59C60GgM//alZbvk/
WrIodlcY/taHJbR9OHq+CTzlDz/3dOyjduKzjpQHDwUECW6PQIpBftaK9kdU3YrmrvN7KKWHKCNg
Yk3GTaBcPlghKrt2SJeiRkgrSO4QEH6fYyAPlunDLrzc4+5AGh7shmqvLfRKeJywiOALb6g5Pba1
gPAC9S8b7zoCvgUWlftb8fWRBbD0X1XsA6ChmzCRMKTa+1ZqKaFovdoS//9EWlzEFMVWbmbdXNeZ
xBm77AevjFBNQQgJhNUIg+LTKxlPHlp7HFBgoaWZV33bYie8yfCj/aLc3Zd5W4l6ZaH6ozQvk5e3
I+zFOKUOIoQc3DLxPQ3Q8Gol/q8fYzg3Bq5WBXLWu2/81XOLsn0db9l9NVxyovVE3SZ2SHOmuypi
Ctmujor1MEDRI0dV70+HR/hGX2TKxHCZNvcTXWjjf8wOsAXfnXiYemSxxZ5qdR7whJEs3pQjwdSH
VtnVXvNpFsoS9p+8XSxaCGpzL6IMxBYBot7BWQzOHZrAxynA80JFw4av/qonGsYYftCjmHkjjFZc
UqoL1fM6Wpzg8OBCyGel4rYQ0trn48M/rwcpdrwOwTgsU5C4MKNzHNKRSKhL5ASOjlLgFHC+7TE6
3oGuKn1HgEpmkQajQbpuf9R/oM99N0tEbIEHDm7+si2RnuP0RRwgd1lxOt+PBDYUpKc9Bgkde9T+
ccBtgSuhhM6j8+950qQZbVf3xROO9p7xnDfV89VgAP77J3OvOY5GEwAEhN77fwfNQp52aHence/Y
/v20If6AGb6XAwzkCcdjUnEkO5MAQYlIj5IMP1RvAFi6xU44ta2Qjof5KbTwUr2rEV8IyR3bD6ip
EXXvGmvAhzjsK1dC9jKnToSRmRHaV3tMMkEXztUSuJ8hFyDv+yVPi/JsGYBU59IWPTE5nJAZXULc
49mS3ZoDlCn5OZ9tqVRKRTweRZPagAmZao2jf7IzQFN2oYZoGPMwJNWx5UW8xSRZRAJuEvidKy/O
oKI/8dQ0SX2JigdLociILKoDpLC10do4PhzigUdpuvP8iP7Sb0HjmUF2pgQ1nqpr7ZEvmyvGmXuy
hSiWFqB/ehkKofJE6l31kSLOLe0T4v/zT92pCjSMwySUpxo/qZSDv2QXIST/6/uYik8KI4qIdNdW
ERgO0ht8orxntHnASJ7UmSRMqfeGbR3LkAF4/mwhEbkOP6TawutcGfFlcLdsuoik6nVAJf2kPoXp
OXuSpKCgWh0KWmVJlZWrsqCIRFJINmpD6AAiCznD1BSQe4twRRgz7rPMuvWPFwXn7/sW4A+88MfP
/6ow73BwXDKtPFQuFyHbb54r5U3jBWrux6ekOtfwr8hch5SnfiOiPFCfEs2k4Y3y+qFqALHF4WbQ
ORNNdK0mnsHbrxPHENpfiv6h+FshMTwwynI3Irrw5f8ISx/grUJHpOHHoSEVrXiMFIB8Isc+YDHZ
5Lr8vlwRD4IPkQs/w884EMgu60NysdIRGOakHVdqKAj8j59hn/XvlKSbn6Jksl67WU5ndZOCi2cd
C1HPf/+3SN5vxhnJqIJjmtmuTO2cpsCIr4KFOctyKq8fJuyOlTiSln2mEeP98y5EIKbkaLgjArH6
jF0nVQ6C+y1GhCauR1TaR8izIYaLSD+YOsewe2HhaAH4j7crVWlDM5RxUZMNTGI8jToDhQaoPIL5
ZCKSgHRerleEKKx3Q1l+jFhhsmML0b96p/yj3NWupgaQ/IpuQkCLqmARVvKKZx5CP/wgCGEsjDOd
emnnawIyNgQzO/Nh/AN3xZKelEIv2RpZdBrXVwLrsYTw8Tp7J9zmjKXnp2o0Q6CtQPln6vnQlYZD
xyv2ohdF27R2oPnQgTM926HVSV3wIOKTNakyoPfwlV6iMUxzhPaaJqX+H1pbAn5T5Hfvqkvc7cmP
6kIL3nsZkBYlID1bsmLtyvsFS7PQZipWniEcXGnb0G45Q5HhktUhUKjG5yAa7wXACp9L4KBur3Rn
Mck+Ve2fFhJg0nlOTK35MbLZ1BQVVbCPd8HS6x4gIosjzuBPHWuHk4CSF+Qqy2Zmods6YUvaysPh
7OGqEhw7QqUqmpOTulg6Akyltxk2uZ2GZrdvmQgjhKpu+MqxN0E50djZ2EysVS9gl5bxBhud2XEe
OAYLIaFzWIO6PKvrB3k0aSc96Yj6h1JQlIoxnDUujUmCyGeCBZuEakwQRuwCOed451FPcVY7e7wY
Pntgy+lkr9qzsl6D7VwMf8b8CS/52Tnlviqu6yxk5LZZk3L6hSDgsvhruG5OhCLaXs9ll5G+9N0/
75fNmqPy0WsKkd6iqBVMWigbtN48/Z1aacltz8vzR6EPx047Vf3uw1F1X9dlRWvKm3tzDLmq4qqt
V61Lz/jCEqIOi0ZlfbyMe8SoRXeWCM2S9CPTNaIoMSUuF1uoDUAVDUF7HNcgp+tVd6FrqXoPJXJq
PFw1/zOffcv/paP2MXduDwM+L5JgNc7FnR0EDgur/XuXv9rVJPkTquJ+40UxmEi9wlSWy3CkjFAa
UYI7eocHIaG5wM9igB3J9juuIkCdiPe9Q5hm6noiXJDTh1PxCM1lPGjwYVy88HTIQM/zk5C251Vo
xxEEdvY4dNaEsqVR6EwaQ31rEjYl0Rr7Ty8PIdQ7XEiDTjP7xyZ3Q5KaE6hmpcS9bW6IDqORaPJI
8eyfFOY7GRV2DwhDsT9mcissgaAqSt7uHtl5ZSGDjrbUPJlh7hEb3GmMFPHdX+3dR8ENyRiWIJbn
1mmrWnGkvu67zhiyfU1ee+VdcrJNsJD9h5itHNgJL2tYEgLYL2/j+ApPkC/YUX+ozVTK+2QKm2Zx
lz+TeKe6H9S8I8g3ad0QG5d36UPo9fhpGMzS55IZhwdmwr6K0vkvmzmZQ58bNp6Yd3JUkMOwr5mP
a36dzljmXmOOxnd1RAI9lLBTJBtOknpCCYOAVVAZ7gGIXGy/rQiVVEsOytIhhKrAbKcIWuhRAGHw
vor2ThN9/nOXWK1dhUcbFw4ikphvi4VFh7Lzl6Cpv0Lrcs16ZeOVEzIyebQzpFAk2yRzHvCvOS0X
O4Z+MUxb/ecfLFjXIalwsl5cAMg8wIRc+U23ySsbxED+5esUy/1IuKWnKLWwaLz45qEwOUGdLlst
qx298f9tlEO5qmGigxsVY6QwKBR+9h7oDXw9DsKO8YC1cGG0ozAGnP7WRch5xDmrh4HWL8Oirnc2
rEFMmfC+zY/suGb65/34rerJR9v3N4pM6yHTmnJpcuIiaoNdGTcWaRv9XFKHnmDSx9rbDjiMQF5x
GUEFy/o+e2zYms5dFrCRvypYUObfu8+dY9/ohcw+jsJswp6JS2R3+9l4x99t3THBXVkDKiHTjAYw
3yuVJMHq3+0uG2H3JpGgoHhp0zvi3EiXy0X0Vea+RwBonzsVE8fqrPnmWE8zpOtdIUaTavKWDeaW
OYHDZa9kTEfqF0m9p/++Fm3c5ayeKY//13xT2QUn4OGUQHnUdLshKHQd4oU4DftWFYnwTNdf5iEC
ygapHnJcaLWx9k2aEdBGf/AYsHOzVYd9vaak4x2LYHdKfGmySjUuR6OT59QD2oy1P14dY3CH4oEF
fMaOp2hZuXQwZ5nBAOFH5FLsa4EFlXfNXbvhhP51DfHGx2EYZIJGeicpS1YZ377QmCtMbpIEaReX
oTrJkLBhCe2vRuERLJPnTGu62hqRs/1f81v0W63S7EHZ//N+DCDYnyzdiT4K8MS8gsSn8Y+wzPYu
231y34lLQMft5pYTzLy7BmpWbhiYPgCym2ta6F9WHXG/ZRlG7Oz4P8IPgTo5oXjVMto73poqta7S
u9u9k+qivzYx5csbtXu+YDtppBXsR0cf2CUS0ZgB2gCrur1QThbYNpAXCZ+fgZisaDcu2ELggNH9
iJ50YidAkBCUElretgl2rjZa3bJTwbEWMs7UJRYh25erxQEsFodMnW16qlZ0/MejNyhf+HkBVgWp
pndx8sgJ2Ta0NUf9wLhcbias5O7cozl8bUSBkCgatf/8fPiRbxHWmfjjuCDjS3tyJAckdmOOErSI
FmKqcLKSXJa3Cwf+TFm9y5vH/rNjAge62j3pTiizNRQTQls+dHUTUOmz+G5b5qMjxquTDNEwvXh3
R4noXlS7pQWpXOg9e4OlmqPq4RZ5o0aEr44e4L+HIr20mQLU5m1FdThW48N4/BcPzRoLif/bGTvC
jsEyFLHacYb74Xkff/ZCwk5AXMG5Za7vus0cI6enJk+d3rJus01OcUBaYa6Ew3eN9EhWfmQcTkbj
ATbY5H+gI3ve1RuBxw4netrPkj+h2Dwtgtz4tvqigFf7MkWRkvqyb9PChtKCP7l6UQBXgA0/ZO0N
QBC0ItDauFdZUVdGX4/ByfHBOrUqI2l8b28CR1DQlcrsM+MhdjJ6GHCW96PlZpEdUG7rNoLsfwNz
ofRFo9VylDh/A5NK8jQz5U6ZrX2ymdt/dR3HbHGluTAdZJNUdYE2sBGz2NCPV8Eyfv4dUv1LooK/
6qzuJaYjio9m75mOSguJNCjtfsfMsUO3ykEMysZaxqoTXcwtMqnGzZ1pmvFXMnL23UxHtps/bCnJ
kcu3thYsFVisX2amgBr9N1MVCLPjo4SutubfTBxyfIWnFGz0VARt3+IXp2xx3Xc6Pijf52RZyhhL
cjW36PzVVeoyjD/xBpG2oBFfXW4RR15tWjMlATv2rV/5P0FUMLQrBgEr6SBjITdF0L3d6A9Q/Ann
bkjQXTx/znBStBqufuDDwh6On91Rw4u3KQIKFG/JRCHdkbJByH2fcOoNpUJOHnerli+pOLjz5vWV
h3SGL6KgSEKJ5mquKEurYyf90Zxsp3QXdVHteQxH8VS6uX86ZG7Liy/hw6M6Faed1OAmlCc8wxvN
/TFo75op/N8rpLv5pImiG9S+spYVfn8t6/HrIdSbtsSVxW8jWHFa5eDxRe2AHfRBhoC9yCz0loc/
4K57VA7+vaI5WjxPPUs+zNx97W20oOHMzq6TnzzYnh06LKZhR5+3N7naTubodYATzN3FT1ppgear
mBOkGjNyq/bwdfVl7sm+402EkTpEfo1iE4vpUNRyd1iDnCswetM90oklltzOfsq894m0SlDbjEJQ
ONOoSuzmbXTZS6xAPE/2gtR0U66ju2+T7bxwTNTAGia/WsFK7MMHJPfd2Y5zlUdywxUNgAsJb1zx
irLh+DbXjS0+o3WKg0KtyLz+lEyZ5F7eepfCst0UXdjYcNM1k7bdKBE34Wj10VxXxZeWTJdqmsjT
iV/gnppU1+sciabnPF63S2fdTMaBtV5032tpUhI2X77qzpn3jpSZzIp1RH5yKRbCvbRNF3qEmmvM
Ot3lfOLfRXt15QWqX2J0xpl5Q+Gd1ohaRblnsoV+Yyc3YJeTlQAnZlNQhvkqXYPBfpIJ31w4w2jX
4PnabD2+JCN3kUqizp16riSbbP2yVghChZz1Ykn4sjDuoDMwuLMAxwHRNcbtb4vzJMLFsobIU6Uu
0GRS2G60NMJ2MNJ3dpniaydWMbhS56cxmiSX2Vqgg8VaBXue/iJjR7Xxyagw4V/esSSzxrTa3sjL
bjUVb35bEq8Ggi6B/TV0iAXSAb0bHqAmvsXaZpgW8nJ8HpqKCF8tgCzwZ+ctG5i8XJ/ecclh4wKb
kc2VUNZF2pO+/BONKx4Sc5GmQa0xNDAcw+crONl8RRQqibLyq5qENqLDG3j3lbEubypExyvr1JnK
fxHB4QYVVki+3TUXmJjoiWxFFGycBDkJfdIHZY4I47TUGtxa0KiIv32KrekZeqKSF2F/HwXJfO3f
O2yrr+KGAFM3rqJiEx4pEHg0Gj6IoML0M8jt8leOvPXfe7GEJEtghO7lsWZazXO1JCYv6ToQJb7g
IED/sB8JnObMsIfCkAFl2nKbeh8xUlpBGh7zlSdTee2B5cih6viJK403/dlbOxk+vEuJTZcxBRnV
9sVN7FN4SEfAV+Dg4sDdartKbZ+GdaIvqlEbHNj7Mn4DWuwniv3ImXC7F1Vf2fKbcMMhnoIDLbIH
a86wd3oWZ7zJ4UEXGgVTKKfUv6trwYRIFwoOZ3zcDqxPGoPeIp6rI5VnRkwO/rQU3l3TOr8zRUhj
yxaadLK8IuP6ZrQ5/xBLO941JqTPVytetR5uouf/m1d4ds+MEdWCFwmzCmffOYJwhhRucvCsYUse
XsU19g7XE6mMTNrzpL9Dye2i4DSBPC15cf0jtGACEMajwReAo38LOHGqJpKST0PJMTlvrWy1UO4p
kPFzQy1+Wi4DDvPe8cCko21lHojqy3/uYDc7Ayu37KOnbKZrt4JSiLPTLCplEY0Q86v0TPXiX5oJ
ADmkGKgegb4yAtCiCVUSduEDzX7Wa/rC4UlgIOG8fjd5bOBJjWvvmOX34fDTkoAvNGxPkBMnmYO+
bwYeQRQXQ96Sq8q2GZKHxHwoyXa1PaWp/c/v4wNMd34rV3IwKWiXcKchSDbqBtw1z7ttLKvdJOHP
5ysRm1cHQg+1U5WqA2+gPO4QYwrQzCQNQxMnST9by9t1KB8gYiuQjQgq8+Vdeosi+qNmvUvhGOa7
cYz5KBTkLDn6rnADeVZRDCzEWYUSgah/AAq5Vf0OQjU1oEBb3ZZAFJDjBeR9H1X4USkcV/vAyopZ
BxM4dQzdYbAtN9FMgDgO7YIxAVSRs2upMxsxloF39fy2AHTawd5UrdbPWjT6lhFaeUmiKmi0mwZe
UMIg2y16+qag9Pm87N3AF+HieJO6QcX7o7ta0NQR+N8ikEhC/ui53wVXKXHiDVWZfQuZH4MBJK92
qRqceKtBxQtqtPptH2l8TOAtOAEmJNPdM4Yrea7Gv9q2l3E6rIervQOlaq9aNzjx1Jd5uO6xzBzg
Obx/4+/ctllln/6jOYnK5yGNt62EHnpfGaryLP62Q9wgSuntinN/UUYd+wXoBcD6MMuhPpNT/SRP
CMj241QsOLXoZxgfSZ+0q1XwwwhzG/6xZpDpTSAUNo9BA7N97H4R03A/y6NQbSbbtsYAlWd7olQF
AslYG4fxSKr5ePAGr2rniZtRpCK3zSeVfR+4awDuA8JAWfvBqDBNQegzoc2rfAUJmsq0lafHwWuC
Y2IsULZxs4kWTpRSzhjQo97ceNQH/iCB9pSYasp2PUrzdEM62M/kUUAitIF4F43DIHNSv8bs1j25
4U6vAFDlQYDDCEqTTqDyWe4afYGZX8DpODnCTPaOXU0V+24lidsnYkGAXKTpwXtLBZSoSq0DF7JQ
iaGJNPvKMiXnaEydYI6Jaxqc9Z3gEq+0NWIb0nVK6n35Sq4lSSETl9H+BY0U6f6+xiPFOVXlyZ07
oEvFRwaXNJMz/M2Jo+Sq9/bxDYlgnay2pST3TW/A+DqwNhmTO2dvZEAP43wz95oRW9NHzzAcIdeY
3tTBj6hJ4G1/N80CZfJff9w8Snvg6V8CHViFjLxwgLLO5++L1pWGLz+cPS2ZY4sOS8i1vTqne96q
//bkcI3stIud9swLMrav9eIrUz/gL0MVmP2ueCe9fNEnldpf+TX1kiqW8rmjgenR2uARb1lTjCqS
Whpg7TZK/byO8qIqwCwbDkFOKd0/7+GtfCVyYqea+wBkJtwm1Nhh1d3nN/qRbbHA3eX5kRkIUW21
auoKAVBAttpLYxhtkK7pwG5RLvOKnesFhi5CgiXQtnUnZxtESXBBM+lB0dtWHVMcq3ox9Xz1ovhs
f5KqrjcTEJcB1KQ9Qvqcac6G3O9X5hdRt02J995INXCyMoNHr6TBIlo0j0oCIPsyfr2jms6tt2XN
PIAJTw1qf9YoV4or5JX3H0ruwcTj/MXTLKAlwUyFSPpM78AVQN/MmQ+9SCuLBwcuUFL4x79QLIha
aOrtUTF8Ypr/PcrdaG3BjPnNkRnVPAVL6eRYjYWy6NNgtJ9rnKD7gb89xUqVqcIhizVP5WVFQ/lo
M8QYqtkitPoHPvDGzOcL3OUBWlyJym99NrWRlHxLHGeZZBvMxBkn6sUS17juIvx5Z8et7YOz4lN0
o+EMVTI8tdx0q+bryKW3ypNDmUgzVO9AXuyNisg5g5Pp0soY2Xt35d+jtABWnt9OGYhx/JVV3I7O
ObTuzfjB4zXInXwnsyiRGN7+vpFfv35ahKfJUfesCp5+P0r5okFHiPyQXuC+gO5i+345Vl2a8vPF
qLluDnv6X4wD9D18bmvpXOU0yALOXSqMnj3d0Sh69LmVOygFsF3XVy86UNAOUz/2E66jmYTnlzbN
WrDx4+IDycyHid5Liqq4fU/jra9nJn+6fSt4TyiA0ylEF5ZgylX+2a7hjG1tAoIZCXoX2hfv8Xwm
r5mhw+e2MYvAhWgVg+gycvWw3OdMv0zY0rCm/pzkvB2QOvfgjuwMJKImJJELtvQMs8mqP6QS/oTS
JXX1+OxnVrWJooqHOARsi1ohuYOHGkAcWlTesb8RF1YdaoYH1r09dxOWvgzp1tnLq8kj8ocYdvNw
wYKDPU1AE96NpKvYLA4AVwqWE8xo+2iiMhpddi5eXNjD43DkdTQsHG0+IOjzBClQxk8fy1G06PcQ
DxDIffeRRHCG98p7PjeZcb4rbFFjRH8FLcZcQospBeOxSnDRiyP+h2WWhyty2lyiZCYMi0UM3APP
SpDdTDZM3E8BvkVk1WnHGkZG/keUsyfndluYS/DFfm37EKMHPnb7oDlgWBwMPlvfrMV+I7/mJCbK
X315Yn57wvbV/e+Ocy4aHeROuW/8GgtwtaSJuR7VNx7hkwJRAePA7O6DB1KIdZi3BXzwKrwmF/l0
LFpN9Z3gYwQr/wIsumcCotvNfW1zWkjJ2vlGgVdK0qKOWcSqY/twGuFmJ34mBNdVu/QjZrp6JSKK
B4wA7G4cPHZ9kpLucEHOPEP/VJxJHhnFf9noGvmL2eZatWERJP5i8dSwXsU3ORzDsZvjSihgq2kX
HyWb/6lhXShQLC69clZH10kpEm8hpArjjvaty82U9OzYryf0vNCcvUU/aB9eBKsbsCskYjSrl0tA
q4GYE7wmtjPFikL+GSvrjhyO4fbSg+CGLFiA71pTFY39oxUU65GGxQmRA7Fa9RF5uoSUDOcLUEf8
qg3FUN27fS0QDkr2wLyOwI0LES9ec3uO0u0tnAllJsQrg4rC9UM7j8MGGj2SZ2Fjua9pEE6zZn19
ZZQtDzZEWg2fwPsK+GO5IHJDBenTPpVgdrXEbl8DUvAgngurSCAQPQuFEorUrkzY3CB+wK2aoxih
wCr8OgxfW4MbeRKD+Vfa3rY3VgC+tsXnZIIEQ9Sp+BuBfd3xH6fJ7ELAUFpGZi0+SHe+p+xA1N0h
gGWfzPHJPNiYlwfkkbZvUF0+VJAj3vH7OxT1BPFTSZLEYqbdg5jPVLd+zlkDPSYnwFCw5zZssz/2
EbBehy/f0BMJ6+73uHd+olBW67zSwnheq9BwsK6MJ00zq1u8xkCXPuEb/heMVNNCR7xQCE6a0fWY
3+pZxB+2mW7mAMR+8deSQGsvrdAywSjl7TeznPR89hv0VBKfBxnhnN178KjUHbokW1gm+9bq3IZK
6WGUsvFvf/Xcgjl7SA6qPy0liu+i1n/z1CWC2zliCNvX1of2xoda0RY/N60sRCxSbAMDqEhuuMOd
vC3+4w2/xxglZdxvetvTfK5G38NX21yjSFyX/N9KxKYDbaIrO6fApzTqYmN27emUZYLzU3hczvEl
CjuOcO6kwbrj/iaiI/HKPN+PcqutgY0pPOsOnhfxDk/tBS3hnlPwL2ohP4k5RYHePSaQpKOYB7Id
ptCq0eYlimUtuB5AzGu0Q5IuTebZYSM3KvsuBhxdCdsWpFhhB/9bnO7QrGPhWnh5judstqOHpdCp
DPqmgQJo4BPJ/Xz0T2fFywFKgxaqUGE9puXdxn/3uMQ0MBFfC722Dih4uWVb3Acj4i/ezAFVg6oB
MK2ETNSFi2HWOJwhYE316F8KMtgwsR6Zi1WQpkhLPhYBiK8v2ti7SxqT0wEUvlEmbGBueieJzXAs
SqCyeCx5CAO8WbZqUjighbEhOoOw3UVerRGWBONt7p1Rmne33ddYMQ/kPyjHPAu5oDe7BrhAspAU
o2zMN1SUUXDBLr+d5i29aVcsJ3Rz9JtCNG64o/ACYV/ABKTDtK39/zCgaQLYLwYFfMzFsRyjwEkg
RrgpuiXWYZN0Dyr02E4m9u3JDFoxT5x/Lzbk5HQov3gYW8WWPaJVZ/83zCaalNYQ9DQGJ6Tskbvt
8cLfoDeCNMOs5SagioFk6GXS4/GywohMfmnpAARz6l+FcI8+vv0bDZ38jb6Q8YdpZeiy3ZduQAYY
o+jch4Hh/t5FPowNXXgUgbw1SbhiSu6VcUBo6n0vSMhiPpf29y71RkkiiK6jwWxKpnyW9pL724wa
wTxv7jO5GRdg+sRdXO61/dmvUAeXmeNIl1sZtcZZSCM5kepMb4fOctAW+nVrxW7phiaH37RhJIIo
c6yCt/M48EvNi3v8WQwSzN17OyYAK+ujEkCM1hry+KgvICivYFNtWzqswCFAtYEuXRLxyOVysESY
SezEuVMtcEwXsmqfzrdZ1aAu2Y4VWkwFtmAYKNHxZUJ7DycK9CLXNAkv6S5tEJYAImK0At2dI2+n
HTvgtXf4IWBZLPd5igPW+8s3RC6DnJElSqbDGu1//VQjaS1GQg9OeyhZv3qvwDd05lcz3ydD3khg
MJClqnkUIbhrT6U9VsSV/4gtevhelNLWiN25yUbUhKxdB1hTtlcg27ZieDJfiPZDULyUgoUBKVyB
8VtCekLAciFvSTqk4fNyUN+rafGuWmAeBibymLV6REGXIoW/IVdNmxOaPjAMtzSfETtTBvUo1JLP
ggchGL5/G5H50uCNopNCy+3vnF9iFM+3LlQrodK4YEpMNvWsp1cydX8ZHA5YAfQmuMwlbiWNkFxE
MTgcSSIH/Mt6VxIpJWltbC+Q7Dn8HtRed5dbrUewbrpSLlASe5zQsOXrkK11n9ttvYky4s5ZK72V
guu6S7gN5QZ+N3zMm7HdkNpaSXFVeQwlWMTDpOwrTjkbcpvYhrHTDjweXsK4/Q5rlSnS3KhNJVFW
B2/CIMIc+qV4gYW1nmIupIt+B9NLhrX1CCKN49T/p/NtHbUlH5zRzJd6JDgXpfNcCWVAcK91YDpc
zM7I2ZMeNeid1qdydwURcnDbiF8fwt282HFDUGmKYYhu9SK/Fm/31Ms5WJft9ESQaPdQCEre9+jj
OGgwhx2WPLlLDD1AHLI0wUWpT12tyruHtJIFNzYUsdP15CU/btOhfzUx2ztGb56y6DEPDbvR1Xhg
W0blGX6PfrXmO6uQDKcCloiJRrHCXOw+0Acg6iin1LzQda4UXJcR6OB23OIdVJJdvBiX9thk8Efd
m+RpDTnNQf0QBvLRXfcgxkkYIG39DUxOIzv27FLG75JVbKaIz3jfL6On0936qMC9WJMSXF6WbjTN
ennoZhvFnCuCBKhN3Vy3rg70MnFWv9QvpQTWIRESiez+AcmOKDqgdLATPYuVCDY5Qe9AERuM2awN
Fbjvxdi3BmyivFZstkooXsWwZpXQtNabHdVdt9h7kHx4gjX8sbrGd7ZjVDNdAQrs+1dGwKQoLnn0
Y8RcMVFjHKjmn3s9+G8bSr+jhJGkNAY4uNstjxs4jOOzU8ibl5jAUtGneF2poqsADhV0ZJIpHelm
EQuvvHXzX1NEzqVNQiE0jPt3Xg+EPg8PhU+m1poEzTe/gXp39UQnoBrdj0IPuP7VDuuhVAbElpys
PF9ByvXjaZoDN9PBeSDFVZ0MLbxhD+xKRUyjO6DvTQHZ5YCLQvSAZUkQmr48O5Coy2K5OwG3N1oQ
5S4LmrwofXL+D+XYEx7Dj/EO3BbtuishW3Xp5xIyrzeyziyFqF9m8DTFX9cgincGeAOsZFSpAhd9
aU3EgYmsWYH2GG1wnmAtD6LKbCe1MU0R/9+8I4wVpAlTEoxLqtYakmuG7IPv9hbfnbSbXzgiOqQV
JOdfoC2Iq18qYt8A/SSuvDNEPW6TbyYrkRY3K9h3ioYDOhQEbCBjzf3223OWXPIGUqTaGrKPE8UX
NMtceqdvkcLUpqlw2M36PDiPWlqtO1/9Ik36y0FH3FvYIVFU4CWB4/yPxwV1rAgqIA4cMASqMFmB
UGmOqxAh6QOjYcflo21Erxmz/L885hleZ2YZ6FHZr7yLXZWPnIctPuslMKIW6/eP/Pks2mUurgeE
0B7vwp7H/G6kbZ7DJ24Nyar+n90QTcLLOOhElZ20SSYbLWRad6AROTyiFpZhXL5hOX3xiZkQi1iP
17j/Q3qf9BSv8caQ4qm7eegu4R5qwN4lushDLbAHRrYe4l83Fwi9Tp6rWQQtemRnZepCt87XygRa
XC88bk1dQDfkMI03AeneE60A98U8a0/r/kmAyUPNwrA6TBwcJhsEvbsMW4PSOjt4Quab2qKnvgfA
csKCcC2Kt3cKgvx85b79YUPE2ebkJ54kt1C39H5Lcp4dogFJxAJXnjP07NZ8lZujkMs8+qqkUSbS
Zip2ZNK2m5HeFoaCoX08JXWnP1l6qULZvWkl7Tfiv49ckF3/QFV816rKZHs2F4NUwyG7sTrRGkCj
g9lh+ZmcFBw7WOB6JIoasJQvcOgcNQciJlPT2vWBNm09TJlfexwRbzcr5NlxA9JSK3O/UXJZvfDQ
F4R/G+g8XsWN1zNtUxxuA3kgB23d4ZWIHgfdJhtWTg8r0b4yj7gfjY/oEtnNJJ2T5Sf4J2oL8rz1
MF8KDwVm3jIaeffzAxs5nRe7i62wV1BhXwSXx30w+T/5j4S8lE7fWZQ86U+r6oXerIkUTBUD7iSq
hSHdSaGoz2XGRpgZwhx8DoAntH1ktopeeIK1vcfMxyGEkcAcQe4XTafVG3K050tePYUMxUAP49E1
D8GCR2SUkCGsl6VY6j2Q/ZaoYB7Ru5+YP10Q8NQl117XI3/If0TPipSoeK9QWu7C/+VKewphyccX
n5L6ShRDGsRzxWYsk7NhvKgxHey2VlPvilsEG5I4cySvJZLsrxjQ/wuI9kjkdm12MJGHDXzdBpKJ
pYDcjte8ssDgT58BdwHWytidhUC75pT9JKU1OHW18yZet7xO5ORGRxKuCXfCiAKmeFzsYkAFlKiR
Df0kedIVvFS+P3/TuD8c2JlbGcBhUas/gyB1j1doPA4IKhLWsknSUgiYnGHRJOWjoucXy93c+2YO
M39RS7S57dlPW11qFFBfxKcy9iMSP9e+jWPSQtWsln4VjM0aovGRSdmACQZPjBVJBKGFdC3AQlY+
3rbNqmhHlOzo90dih3WISDFjfAFvGvxJ3CPolVKqTYjFK0QbdWtTjp1BjlYqMCIlXnfSIGsv420s
JHf7bTXolHNjtDcyrN8xnS4Pfyofd/MM83hHSL2xkYjZTo9LzA+qx9+09Dj/2Eie90wDv76N6bDQ
STkbR23mdLiB05cM35Wrh2GQWZdkqCBkE29ZvP3vqVWoZGEI5FM+PJfhNTlS7D7gVq17LHoj+zXA
KZu7MPLShcsIR2jlpfH6LaY6n+To2yD3h1hu/5VAL3mhqB0WtPGHcHsqXW4ZTMagioSyuhCBz29v
54jW58cYeANYpfQK0RkTyR3qaZyvQ4OGd0VulGGgVmYBxey5hmgCWxFqvYZQJ0e/eMdNbhyDoijK
TsKNQZoermvka0L2MHLLdviJBFTp1aVwGnkGu31wkPcEovdv2O0Av2hfIXatWgrE0JAu8eo5nIi/
BOtpYh1asypLEK5aGyueW0bXZoNc/h2ghvvMWWoLftU42r7giHTkrUePe3+D4WILyeeolWM7QMpY
13kzzz2u7AcDy6jFB1Y3ODb4sOnZ3lT25vPWAka/Y9Id4TheNqzskqesdMjNZk6l6Hjl4BsMPDEu
4Rhg+5S1jiyiEBb9rc3oaoDx6NQmeSDvAm+lj+w27Ag4CKy3Usdj97qKMuNSA6nKgJ5w+RkmV8sR
GpS62hRSgg7r5y60DDA9XsqEVrhFmGV1K14tkHUPA97KcKzRh6+b5ac1H24ownV0al3pZ46LUjKT
fp4zJAIIYIpFJzD93p0pR24fuKucwx50cCN19xMjdNjJAWVp0DuuXCRJdTzdsQ2uxze1yxtCjN5p
lRfQDi9QKPbMP/7L8OEiQmxLlmx4zuQB4GDpRhGoMXdoWJcUojCzrfkPiEGLsRVLtLlWfboZURte
PzqtCbM2R4UjNXC5TC1SNFqQkfn/Nc1vKBAOTUmgaB1Vbb6WXDxlW8kuoikhrxCKeZjSrW4p0rLg
Zxvc6gLDvrPw9036UX7NJdndGu9FqV+fqfKoKFBbWs8vhvCGVbmZF8bc3vFyJYolQIrS5gTW1yBZ
tqHFdlWtMXIFtXUw5krAO/LiaqRBuDH8NzKK54bB+7WjOnoWM0JQOanTQ5D9aN6o9nkCpXbMrADL
3FMY/7Pwfb2+8q7/NE5TfMAkZ5leGFZ4YR5Qvp2L3NMJdQIrIJkEyh/Pz/PVkqT/KzIejIersY6f
y/u7OQeWKcfFbXpIeQYKmi6PKhFf3Jdp+0JIX2WVOqhRyUOFm+bJwXQu1HDdS+8IWRthl7qA6LH1
iCYkfShZOgmMVxR0xs7Mvb8CXXh5u4JKHGFS1vYj0zgWquvMjuvsq/MwHg/ukdGc7GuGkAlOzSaB
6N6pCwxiqtKeKtYk9NUOvrqXPppxy7TWsbuu+rbex74BWqqIe+HGP8/C1pqlYSqBln9vfCeYKfqq
t3ZeQ6shl9K2xn5SEyMQoasdUX5Qsa60GIFj6U/VYNssyjloWg09grAuw8LRKY2hiUrdrPkh0MRX
6/RJGuvAvrd91f1cTZtXM09wrVvg0nd4vgglbnWE1gdY349oD2ogIs0C1T8KsCbvAd7v4QmC0Sra
BIzkModeqhsxWZ/2yW86mgNrrAeClN2JbcMbcQg4wdw8qLdeWByl+OF+XYtau5vQxOJuUWLpvTTr
qQ50slVKdGcdoyQ0aqND0e6g0u52V09s7yh44LdeScyPx+qjKtRgsf8cC/aSd6FVBHjQ9F1C04Ma
wfNHzqZdSy9vvRuMex5/mWfv0uF1tYpHR/FrwyVE/bWYfThQPQUC9JU7jfzfwBOGRYf3lVodatrk
p+JpD9ufk0qvUNoL/Z8AarE8U/EBWmvJIBZc16QAOrK3d+jcdKOtcIjwPbe47n3tL0pyatlVA4py
CPt4jn0Qkg69JciqvCmiurxy/NrgY2rCP4FfohhVqM4MGOTaA04S6/GnnjERJ9RcF2mhvOPHJTpS
jR/g6DAe++sfCoCfGoYG0tgqEQABjjLUDw1PJ+/PWNDMerFiD6EcHs/KcHXO2Jw3JlUn0XteXVH1
SholFoKq2ilufYJw5TfBnUb2n7OP6aYYYH0F7t+ODCukn3qQlkmFmQeEPj/pPWMhP7rrtaM/feJ9
AOEdH+uvo9cliiPpMp0w92a0qv1OjjMLXkSkgPZ9MHo9eZ48HJ0tx59lWS+PzoJTGxuZj1K4Em/Q
e5BFTqv8KW1hR4qDn0KOJf/pq85lKQSu3hJjcNoNOL1gEww4I+CPXiwmn2ubkGsvVP1k+AhwWWRC
XHoUUFaaLTjk4O3GftKUvben/6wOIzcAn728GZSGUBBgxOPAl3mTyNvY4nO6BTEATmUBYmzIjI8V
8zl0f/ORSCjU5qfh7p8Ealfdc+00UYvZxtsOinl19+Drl7Mnh0rPM/zLa3PXPArg6WfX7ZbXddpi
wxmAC8QVBsODgrFU440lCDUAHo1GQNYOO2Y/4DgKHnsMONimcROss+YpSjXtf3r8MAhagFbdvLB5
ihLZLJAJUWeNhtGc0b4L6N90YxZJaIKA1kYfVCuQgfAjZVhPuK8Z6B72PcRp2Elwmfc1dQSTDLd8
S2FnGnqEQXHDX6/Rg85wrmHdkeHVMFL9Zh4S6+glM1AqzK3L9l/HYnNeBTcJuferYpUvDRuZ1Mpd
jqYOye9JphMMS5i4ZXXt4sxvEJWr1NCXoTFKHqMhsFno05lHKglsl3iPeHQ61bVx+2F77Ty1yJF7
qg8PRAyAjJ64dYItfMRtrz1xc7hmG8YfYb0CDwx37KRv2wYmOEPXjl5zq4PdYn294tYW65C138lA
Wid59Nd6cdYRsm4QFJz1uy8/wUAMtatVZhYOf6jkFxdZoSeH5Y6cxUeQq8KHipxZVKEw9LyZ/Gwy
V0vQvSUyBmxhbYZhWHOk6IfI5mkk8VxpQGgHj8Ekf2VJbG2AU4Jf0gQdYVAaHOaQYcbBJ0kiQJDS
U8dKIW2RKPP5rsBYOwXA9Z3+CoMCwESkOR+sOqRj2sabUcn42RwTKz6qYG7sQ0mN3AzH0orcSrf5
OHnYywpfK5cmN5i8l9oOXOFsUUt6uEa2dGlo//3nq2OpjK8BCBC2JCRo+GoBLDGMEVoxgXDtJzQr
XEbkH0xBz1CtBpZki8bUggt+BMY4JAnKmzmFn3I6atFyZ9wnWINtdlBotfvVX6MEL3OT8PCeQIpV
qLKRg8F6wwum4D5GjrXb6FOW+RSh/118mP0IjfRs9P3OPrqT+A2w/p6q5q/XXHmUTsGeU2r5gYLK
AhphtEN7pTa6ltOWC4Bk75nRVwPMsJn0wS+l9QSw5EGHv2XO7YLkp90tawaM+NZM5WfwGrI6urTc
AgHoTmhStBJJZ2OqkiMUk6VMKuQzRYAybEt3JyK4b4hm4pToA0kr17MYKQvszQjdhr85kZlzKT7V
J1R+Q3c7aCFOKFE2hW5tcXAMEduI/ybHkImeWfLrtAd88LHchSjCpAckSCHIbybRwpOJEYwOSTro
yu83z0ZGAJ3fK5bjVN0axi/rMM8d7JzW7bYWEP43j9OdzWa0LqyiyTNspMvLkV1WRC7TjWBsFwGN
se4owIaOqBaWo0e0hsEvra9uWJh1tPAW5GfDkx8u4MDYiOVWMA883x7ASBcYAGP38LzIRoZZgF6J
6F5N2C1ebo0EuNhyyjNUJ8JauRcaKhvvcu9+o/CDWBeupiwAZ3HiVY9NxDe6G4toSEGPSqiAsjZQ
5jihv/JORdYptwZ8T9Wk4M1255eBBz9jjLTutrI5Ix52fp5AlD98u4eI619ShR1p7ijWGjZcSF6y
wiL5R7U9D2c6kRqGhXq/dzwG2nI1nSKAJOl11ox3EYFqqs5m+CxUvwllYvHEfzkX5GEdFR5qfCBg
xI6QGuX7KFzeKOfD3cjie6XUUgSO0TNRDGSFaNLliqUqZSD/K6SLzH/e8p5TFOIwEdvXAr0aCIz/
DeXv5NDkUAuf39HkFGHZEZSOxFgiiiW8bvpCRahYa4mrYTE3d6HBevvhhRFL7ZT6Gr1j8zJpiR21
JBAgPuBu5DVJw5WLS9tNNZ3DYJwGLH+wVGb7Kf0lFRmKK28bPtduEYzz+5tHHCigRRSDrXbtJXNU
NgCvPcztU4/Uvr8NF2fvSsJ1Fz9OFIoQQQjQUJE5LCKDdr7jxiXtq4bmbZkFOmUfCzo8m0LREFFf
6pjnt3xMGnBEwGxxOkoWm1GJ2gCIOEb2XlAJgUi4CHStf1d8RriC2Es0rG7jbsJd5b+p1j8HdLhI
tsAcKTCLgQVRWnRUM1yzI8V4g8U/EhbqF/8yuoUXo/pRDF4ujM4Nqp42+gwCvw4ZEFBfYCgRtRT/
XrBBDl3WCKW9XptuNDDaF744AO0PykmMTtmQJ0Yky7iE9Ni5G/sJ/9g9vIqWiE/CP8DIN3fO2O+3
T+UnfiumGksyOan9ec5UFtuJIKiOGCJAB0RIsLnKJgHm7twE4ShwvBTyyzdJWmgK6Fq5FuEXg9bY
7KjoAIGVMbbGJ+lntb9xNb5MWb77yaL/Gbh+RC62EQjYvMxaY/uz9DV3M9xuit4TPQWx9rPTqh2/
dd2XFmARoSkTkWe4wq6R8SilKW+VHdnTepIi7PV23FG8NeKdN9p+tutQhG5GJOWIqsymcQrvIZOY
A1ucO+lcswep9Jyd9eETd7IWb565TeJhem/bO/48nqae2fQFqRzW5k3wx8wkwHMQJlEwbCgiO5wo
r1RxppWyGhbtRLuzLupQ9J+SCw/DuRoOwHuHyQenBgZjzdSW1aNIqJmPZIoMLRpThI8hGDlNvgmv
zYd4o1PsYbs72PVj7VhFG9xHqtoVu285vc5gtcOlvDBRIKmPDfCy8E9ViwFRUD/MbYcFqoJi67hX
GSIXXPf2tfURwt++S6zkgUZeAyhqZAbvIJKpzeV6p8/wHDbj2LxtqpZcYQtJAQ6uLiQq91wxjuYa
6vrxY9ojnHo1la5KlSwgl1SLVO5Z33/cJQbM9DMdT1HHG0ZTlt5cO6EgO0QKlOR8AwCTVt70rlWP
oZwYtd91L7vrxUFvgoeaqRDuICBt9COFbUyZcUWWjbhObXv2jxBSB78PdbmzmAj3gxVEgT/970bp
3a2YchGSobDwSdQc52CbPlFdlrFM6qN6b8uZCnCbfqrEFRcM7Xb3dZ2x6zRAPdHtezGPCMxfnTuK
fF/nlu73OlINrCeuPrpS/ycDjNfdsgxE4xW+Mp9zCtyZjLwZUlU83Lb4XlbTfHVkcem8x9rxktRK
KHoy7GzWD9GCLWRPkgCMGFS+mAhJK6FgEuzj8BAzJY5yi+jGOyFCoowGHH3hbB3sPoBKqflIN+jL
lx2cJoPkJVO5mbo2Lh1ylZdOiBZIre6OIPYHHxjqEClkoG1utW6Pol5QKZKg2aSwcdEAuaA5q9d2
IcHfHkLesY45con2uIZZH8fjE8kfZlDl6pqm8i4HRHlPKRx97HqB2HWMZvOmVWTeKvQJemUb5Oqk
nQ0TlkkOB9HlyuW+Z66DQpDTcWdEEfNhq8mbhg4SKxaungyF+sHnqcsUMbbpdS5PC3UsLeGCfmNY
K6Bw/YUHfCDggW+1nUQGYafy/ZDjsd9Fpni+S/33B25HxXY6+O3MmaYZmxOIrySOaYPt2NhnQtUF
NIAL4demLibuFPObh9mcPO+qKJwzOiurT+eGeLrCCwwo9nsm16iaVqC+AskOz3dhQ9fqueGrXirz
6QOs5B/UVE6dTjwiWl82Mp6BCw3SB5fA/HqpyG+X7Oo1Wo6RRMnzlCK5Y7ZFUGrbUPV75QklxYRS
V+YY9cW+OMbmASKtZA6gSUgGf1FoaM9DzWwtTD39SRmEIP34Zn6NgWunOdjotHa4jGFuw0nrwqNQ
WHBET+eQq5SUUJiO64VfSW1cATWkk80Ugx5g/kQ6J4tm+3PrkTD8GU5C3SrgDK/mnOCXE8ioR8DC
KcoMbKDe0EBS8XchBI3YznkgM6ih3vzvCdjKnMHAuZDHJ1rAHQtIHZBQjX93YKnM4NFcaJGrLY7l
2disFVCmrplWpBZaRGMo1MxVHGjC6P/bKB451g/7h8tYXQPsl0cWy/YJ/hD9dMetB+5IuEUKlh2e
fn0DtMp+tM6kVv1xQHWcwEppqgCHpULi+i+tjXtaxsZe5q5VRMJj4Etxqwg+pKsTvFFU7O0nZIOz
6F2bsv7Jlu8xY4eIdb3d1rNvA8D1fJ4c+Du+ltJO9LIyICEH064u5EU5RAc+595f/VxvZwV+RCzz
QHGlGJ1dYm3WJqqtqju+O24lQmsEOW/ZdD9g9lCSxE22jPuYw1hfanwBDxuqr1Mf5qqGYvKzzj6C
NbCll3Mokkv0B7r2Gjo7CVr+O8MHuYMvhvtnytoXnavEbuo293eGpzugnO7V4IgynKdvkTDvlWIs
7mgK2Gv9+3W6LC1MrS9sPXcgixINCmpTdPraMS1oGd6sMJYshhtTtLjNMPfkm2n53tLpKIRA+pnU
aZ5F8E/1oa9T0/bq6VLnSohr7hy9iawOLHopYY7Q5wBkgmRVdtTJrZ+zjmgUS6IS/VO3GRwX+mlJ
HkH5mx6iLVPDK57/GVSUnrCcUtu8DZavpVr+cEaRHVS+fv0fHlUGmwNaLvCBgDhV7c440goHWbX3
lME9TO/LhlKWhlOqoERCb/EQcBzVZayIJz2TmRmc1S+G1T/yFEwmYA8A+92+lyAijpZekK0sVKT5
toJ1J7gc1OjNCciMWv646i7P15KHYHb495LWhKI5H+U0r+SL0upFQF+LCnA6OINNDrlp10WOAFFi
OnTosqj2JKXdItZmlR128jWHJ6a+fGvuKqlcMRgz8ctVEaBQExR7SukaSV/MIDjfF2nIv/yVlICv
S+VOSkk9jh7hdu/b846qXLvjmvtLvRjE61zEbi2ibnjd+ZgS/a+4AMbOY0zyP23d39UoJfec4mL1
EKnkNSJxWQat/H4nglVM1MKN3eI6nYP2V3Io61jkBgRUX9EBsBFrc5lOTrOQx1M1is0LvpItErOi
cbABv3OREtGXwQZ+gJ6otCeKYUFRIYWgnv8mPfDq1o9RdCE2y6gisGUntMXE4ezD7KHbe49KuxrD
9S6W/yvQLMX8RMt/bfv7JTVsBgmXNh7qXzfk6kn9qWKZbSylpYdnrnXW5q+Yht25EfjZCnlkkQT/
xm7k1IBQM6og8oaYmsmygjc3+wucLN4Ldeg8NYYYr0pnup+elVhb+9x061XijxqllJZnwKGpAx4n
CSudSy/JgIUabaCZyqxisUg2oaGMiZEODJfB0w+FtF36k3oReFjZZCiK809VUSHhjVG11t7456Kg
j/R2M2SJtPozIe3WczYDD8+CAozpii+y7t/nq+JCfEGEopfoIv5HupUAWp2EeqfpO6vzScm9ZQYx
fTpr5YD1nVtjX2mjUMtjTpdCfSxDOokKLYUjLmMm5vkZu8UFLbSuz5QzIyRl0qwxRC4bq1/dKHYf
YLv3hHCnPs5nDvlsEdbJfrWrYp1MrmLOKWqv9GH9G8zuqqq6wrNnYjauZyKnWqQ5L0aeTxrVKUNa
vgoywg+0aI+4W096GiFvGe7rVu2ZMXv6x9OWpTOuVn7FOwkyv2/g/r+5QVQ0Z7Ypf7UUXQAEZ/QI
ubrEiweFXNp0X+n9XIp1VveoaPSLy+P5jOIiisp4JbqdQx0X9ZBfKDEtuIOkaw5tIAWhx3Bn3VbT
XFC5DVPIe2nfpZlCpA0S4NkWKqaMg62xkJpnp6f4w4+k4KGquQ9Ux6aQ9m+hBzf1ryr71Z9aTtT3
m4/hOJQ7lhzPCJHtqLM430Fx/hDDBbzEeBG6lGRTyPkJzSNhcjF/5oJdiaTET7L/kodOzWlDHap5
0zxJPoVqpMs387nCBxyI0el0Rixryt2Smco4Uc8HiiHgvTWAiHZOa5ovSSe2aUFk3bUI0YrgZjR6
QUc5w7Tj3JFXzJq2SkBLMaCd2V8SYfOTPsgbYd+sX+AE0lkZy758gbKgTNOazEbK987L1W0Y2OPp
qcPtMzCgCAp/wD+UTfi18NwMAFtx/RLwrkkfC3dcTgYsds1RdG2BiJT3dcl3RqhgyU+S9Tx7O60g
ip747WdWoxNwnt1FMzFyaqBrwqS3bRZ00TyLay3J5xmgLnspauh9mcHjWiR3oW2AffmSFSS9nDFI
n+IB7t+X35hnayaSKGnDRh/GgJvXf3621VyObjVhUVgUAq68LoOnGm7c3+rvsWJEYldn12d/9OwI
G5kCnSTX/ulkz8UZ0ty159K+P4tQZ5rlohUcU1jd6CODk7JrH9arosCYXWNfdsYLoeQHlyIXd7vO
FHUWB5pULgvdmOy5l2WsPw3ragRjq6FB+QcHn79fLx9PzjvMG/rYMDNBYrJgPDy7IqDB7WQn8e21
MzDcve5AycbaJTzcELcACVoL5Db+TQBRXQGhZZmL0h0zbEV3fZX9c7eF/j3A2PINkI5gVy1ATo91
wf6xjhBTTpiLTsoHpICh9f9CnGzIOCFOS5tobMTRFlCMoZ/cDCw7srCNgmjNBeMXdT4kjs16VC40
3gUuzPtiNPW1wRWqbwC2fcp3tPxuTENu6v1jOxukGvjzP1Y/Ky0m0+qglb9mFEpVQ0OcJFjj7R7d
DCWNwiUu6eDHtugnpxoQ84w1nxutzRUURbL6eyELjfhrnOrOyXZ01Qmh/m5Qlr1ZSpirIiHDLiZB
j2mfbm2g2GKianZ2xmiQnJc6Gbs+Ddf0/vCRLjZV9NHb6D27E3sFuycrTZm10UqisBXLmZB+q1Da
URybZbymoimXHwjxwceP4DTKYpa90ofll8K6NebIXxcdLTxvCpdjmcSDjCGT+/4oXd5XMh43k7Xd
vRB9bL6YPnD3mskjpcJDmmAMXqRDivqsoEaOCH9aJav8Q3JZ39rsS8f3EyorC/HcQ/60YDVBP0Fz
yzIdWhRkuYGlO7QP1zoQLcyGoKsfIkBossMwoy25yLPeeU1OfS8D837sew30KNUNLM6ZTWO3oQUB
/+6Fmj5tC7e8O33XBqvK8/tNYno77LsRS69LwBlj1UTGZ3SOMbLpX6REYhxUTP580EUJbK3gu9Uy
CWWNN0H7P06RKVvm/SqAMU03oy1Nbl1Qr5tB5kLpKwVEmkQoWI+1jbtHE4PoudkD3GXwEFXBdIEv
dN93t0HZ+xOoxrv8fyrMG89t+NzzuQOVZnnTDhzw8D2m56weXMS/bYMPj+pRET6xESzuzFtoEkAE
Tc9tKFVgGCs8lK896aU3jR6i+ZCp1mw6mUq3tZZ8IL09YpXVewRpJAwSokemvJZRLSNC1EI6NVgg
Iqyr9Yw2kJdlDv6O4Z/xEFdi+P8QtbeK6ShOzWBUMMleutEQQfzE/CGnSoxcUCu7jbbFM5rJGS5w
qmA5URv6EcFRKE9yYLhRC6xHA3Ivg77fNix6jHWoMMpyiyoQgSub8QRmZqi+k2w8MuZwGXfNtg+E
FecSeIw8LQ9PjijRYwllvJFrwELZjXOw3RDW2CNKwgtfiUhzijWOA1QPBu8pKJi8q0HSscYzB39e
GO/5abB0Q3I8BWnnwugPOki0JPqlpeZA1gYv1Axzl+dID8C3KVgdOsBBJ+TjJWdeHUvKN6tbK5lX
5IIkPmfnP0fZE6Uqgv3lICMfBN6WmR/SPrP/yXmS2Nty6+MwrhQY05wELJY1zTbbp0Mw52/t1XuK
UFZjqFPLYja/imkmRSZVosBmeCKTOxflBu1ExwbZtGLrRGWjhLZDvMxg9R1ciaX/v4WTJtM/V6Tp
0j4au+tSsQKU11Wo63NMh6Y9O1bQa3c7lYLooXPvS1LvJy45LQ2LqyGYRnbRFnGJFsp61jsoRREy
1iGVW9yO1flnElE6nJMPl0eiKYKNrKgQ/stFVnDtS/nRvenVdXdnZePEfi4VVNRL8lWiV5/l7Egi
P/muZElpLnBhHYP7nDKrIZffcv0Sq1ATPc4qzS8Cuh484KdWGIWkkSqaj3QrHPIfzaAzI1yIIpup
cp5LhEAFoR5Xagdyt6BsI1ThAXAxpQbl+HnkoAvYz3RLUe2L4zU2cGq5Rl7k2G4WNyy04cTdKfwa
aa5OxWn21hzHi+r94uAUUKdkj23TyC4eLyOk0/TIL8GR2r6kOhcNUyUvFQp8lweryWYQXUlDWbJq
+3P9deU4fi1VngPjkYJlRtW7+eArjHOBOcM2ZBxBrpDIeTx0nN0PlevGO87wnU0oweA/q6aT3/mL
naQMsHNaasgTtpAjvmrfOdOuHbJXwsOznGmzomF9mhxot/HeOmopgSWUss1wKeqN+TgFY8Zj9WeE
/rSUC5h9wy9te6tztbDSnpZEg15w0TNh5oTKMw186d5mJrdstOFc03CstbibUTZRAv9/cwKvvep6
eXMjgXQPMTYZtYa1Uyq8vbjHqiwx1DvpCY09XtWbwA38A2MM2m6QmWDSPUNPSSwb954ImoxFSNAb
Q2lqCf12tM1i8X7A/FvICCR8axni/nFdwoPI/+2gxLGGNdaqU23QMm0K7PxhYV3pTylOaQS1z1Qc
Gb2Pr/+CjEXjqIhpXjf137J84A4+gk4Gmu6+QxjY54+D98T7tu5Sf04KbFWVhSQi9YnNy//iCyD4
mgdfeY7pPA03/YsL6QHrCj2TO3gcEhuvoKx8KbR6knIl8hCqGR+jgN4l+nIGuqbAKwDx3H2sKxbM
aTgXhyj3nBZM6rlvhOIERsQnVEvembJRO+fIYJUyTi3JRymXK0ozGgBC54irrI5lTWi+oZBfUOjq
b/pfsQwXFf6/9Dg0KY21dAGIg+6ZJ03yRkBadAW4wWXPMa3CmaJgE50cdDzbAk6bMo1xpyhrcjUh
bIDJusGVy894xGYEJtqYFezK99LAo+Sn88haUu4Wr0sb8slfErwAEIUkqYgiR/WXoY7UoDKURoed
rJ13DS4aN7fwLRRZg12vFGTw+zto3WGmoY/gK3R3bkmuSHBt2L2QofmGCQ7c6JBq1pkWrApjxwPA
0f0GpzKzOa+yAgmiEOm6jZ2h7zjgNhDOrUzqwTQSgnoOWB2ND7e5gBIo5ZtJlOY427TG5Z0VRXlH
sQcs7ykQ0AADh6ACJXaQOWIy+f1WTHUyH8z5hNgY+7sOfJ5lU9QapjVbrx0Wp5oWtS5uosCJRanv
dHdHKxN/tNElkC4Jyu9qCN+yUMoxkWr6X/DJgORixxn7n/ZxmgWasph3YWfRNfxEyJ7yyAB8VC3W
rbsvB4oekAMcOqAe5t3K3kJsFnrpB8NLpY+C5T2OPkoeBBTIuP4TRRMy+fMIj5+uRM90zzKvj6r0
PMw5ablzfoMxV+iiDOkl/X529wNJ9d3naP+t9GY7s4oOHDVrBu/v26x1IqsDottYPn7aVHMuSlVY
JxFV+DRcQuk6F/BFkcs08of6yso8HBnYmA+N3ehxDH2z4/TbHAhv5+0LP6ziTCQN6S/kqEDf+m2z
UakNr/YmIVG9/jKwcApVfhR74ntpYgjqn/ERXlvJ342msXhYsbA474QFCMMlJdED/p8Wx+1RXjtq
4yCzGZtdFpvArhAQX86QI4+LBCmP9ksqdjjUgQZxuj/R78zbkznbR8qXo3KKymqc8qGs7KcMMlty
3JDj2aYy3JEYWFkjsitObq0wMMKknuRJOwoV7Exd7ISH0dg4Xr1AH/7tLNhZwxfl0ChmS/kb5TFa
jdw8qHvDN/3V6aU3fGOZnyYz3wjfFyc+C0eluv33mNmZNYgdCzMvuxx8FLKjZeXIC5kiWv8bzldI
PXTa9X3pSEbiUw9/cLCnW0vbSRL5GogwlOJn4cXbAZzOLNyy7vPhHNR++giNecFFvaB/CIG8Pnrc
bz7s4ooX9WSFQbLaNwlbMCbe8yoFXcW0uDpGmOg/gWQL6HpUdsCZI8S+/O5ZuCveUbarMKNr2dg+
M4oMpe6q++fjre8kxCU5AI0Jeet4MNgOxCddLJT6rae2qujRIXk8S5viyjDo2mvO1aj/Q292DLRw
vScz4aP21qDHQD6B5OYtL/ZnmjQYVzIgzX9Iu2sS4Tvqh9MXazjr4+e4KGHXnU0VNsiOdcFN3SHW
+hy2E9xuq5CAcI3i2jzPJY9MP4s7ZiNETALV50DoPwd8zH8rNs3LFGjmjLPn/PQtMKyzIkSngMPk
N1gs5Sjy90D8lC2xDs5KEj7ZFQBAe9bh3qHUYjbrahmiREAKFy9o1EGmq4ONhvNWq858lDMAWzcD
XQHqt58K9xLa61JLpWbhssY8iGcf2xCOvSYQ/9QAEi3SweVOyPeDxP1SsLEG1WymCgNv0L1CnA06
GKzbH/YjLHW155lmpMo1h/Od8TQXgq1zgu9Wk5nQ7TR5eF93Q2hPdGHufc043L/gEubs24qC+ABc
hHUTclwM+EOuP4vRpPcROKQKUUHPh+p9f1NDDdIHrrhfdwCh7RnFrQ6pWl9ZGH8JI0vsWHhI8YJf
FceJd1JjAAwgG4FuhQDTAgZho9WojTvM+LHGfyWGStjXXrcqEzOwI1SyHe8nWJ8nvd+3BBD9epPc
52CdzvESieEiyEMvRV/fjilIags4epDjppd2LQLL8cJOvNFd6iBDXUuAHeRYfygFD2eK2WInREkj
8FpUwNffSeeQh/woouPlT5iRulcy6rTbLuSBR6JTUQ159Plxps/Ju3eEfYQkAH1yPbHuOfn0r5lm
uvrs4SvazU4ti3abK5isBiu2GAnE/sxGYk8lpZCO4smjp0kESA9k2VlGxuPfeBOjr7QABms9Uxut
5uY902FPVks22B4IMFFIc9xcDIUqHspPJekjFG/LB/u+z57LoV1FPXDhfT7eP+O75VAubBiOU623
1/PzFbMXPsebx1qKSaOy0Y9o1fhgqHPqsPIQ3TB9Rh/RD6zWmlwtHlPOhqHBe5peXp9WF7KV4DPO
A/KqlTem0UbzKT/1JZsPVYzY5ju9/m9x9YtW7VIZsMcnUg4UbtfPKMXLubc+I9i///Qg+W7eCbY+
5lDUy1570t/l2TX88dkSEKC/SnB6fAdim1ctpUDsng5rFnYjlBkhVTjCoCUGO8v7xczaNZrdIEbh
yYz2dpxctDzhkMUR5MYBalFLcUbTgsG1wWq7OFMNDC285Z7Y4P1HnGIGWq7fhxIB3wT6zM+wvkRV
nknoSBOkglnh/tALrMpu/yfvVKqsm88QkmkYH0e3L241cBHmGtBATc5xoP1jL98q/bsqD7Shbo3r
VilW80JLEjQodD5ZBYCwzMrHms5b6qiv6MWKZ7q0Lh5rcnO8M9vaa0qAxYletR7WFu/XJEHIwIKm
y/fMfrb/bpuT7A8rie6ZxlMmSzsmv1BOERPl3kQQWIF2wuAyVVdxp3Nq+ce/i+7HepMBCzsf8tLm
2FLFpjf3L3SFYnD4WXXpAppJjATqFTvbM4BswUD7WEK9qYOHdID/2CaTIGHYmfaRtYzwVrXJv7C9
a6Zi0yV4Y5YoNGRN9oTy8VzDAJ84+ePKjG/hr5i64wnUk2upgeV8Vq36evt/w2b+vExRG9pTcwev
sGzcNiRSJc/VhA/HWeaLuXhaxSfyXv/Hz4L8L47wxHVLEFHHuyogOYI+TxQSAvXNLpsXkZReGO6u
qufnXoWpjOm06WT/6v0jdI1nm7qToWd83m0r20dGn//FS4A3zv7Rs/9LGzIdKriaTbNBDNWS/Wwr
KpJ0yBarvwxvUYZXz0IC/7xTyO1UtobZPDmVSrnI0Rk4Do0zd8zeqSGdP2FK/pnjwsu3+WJhtF4r
+V2dNfNv38Qr/U7mM0IUIdVUhicFR/+qBbxJhOVDAlq5KBfAQYRSgAQpZpGSSJ+kgY1poK87fMlG
njij5LJDvrHpKlNTZ8ddnXd3ew09Pz9phmX+y4esc5ySD6yoYBMZhD2NhqVDODhNmsBKGG5TgB2d
SOw5tTfwoLWL4ZuXoiF8NW9c6FO5743ax9uchLEdREyO/eIbdYFIV+8VzDyHh1XWqZwfRf7jv6EJ
iUd87anIVSrYL5BvVBjeJH7ruLNQwgsAW2/PEdL45m9wQSZo/45pMfUfMb4pjs/cVNYNYhP7wq0W
JJqMzNuohrOfioGQF+8togfsLTHy+u9bJvbbybI0HUSib0F0577X6ROmfPL8/BMq/BUIy15bw15w
l++yo29FAT9LxWnaApApHcxbdm4mS2XGdLJLB1iICg9GbFr8ReLlNVipwL+COXQtPh7ZMDedyyxw
ThUY/MFWgQZzy8UhwFGUdJ+vb3c/U9wyjf600l0Wg0+0zCQvLEQp6Q9u3gQ+vxe22zryHJo4KZsF
pkzGIzN/24qaGYMwaD4Q4T9vR+dNlee7ioksq/3NFNk6cV+OJknC/Lo+2E94b6LNNmf0gP0YlsWe
lIUB/WfkZTDzAPUmLbvCZ/smXcDgcvYpfMeriaxVX/vRtT88rspM8EoCadkl2MatIJ1RWv/lYwex
MEX2Y0jGXcTWFYp1PATfH4hMxsk0bM45i2D7/5VgZN3Z5XOSBj9x/E4/0OQj8jrpkHJrDx3l054x
0IIbL6u9Ep5/1E3agB6QHS9PIv1tNNTF9rU3UWdev7oZYnD4Vx1zxLY09t66xlDDoR2Xk9r94Eej
o6ThZytJJY9Zotj2clVxmFs0npflSGRXVbupm+uz6BvJEKGQ2NBEdPujOHoHhCXYFR0mAoKePzgw
NS9yn2BaDThMG90/BnL4MamTOkt1HCfeNDuomEimLGRG+MU14OeWcKxPoLqqvTMf1lay0ZiQGVZu
8AyejxfbRQBtDKrCX6/ufpa08n6zoBh2l3V9axMuOjzHkHDC1ZFrxMEzlOh0Et6R8TA55UxkG8hP
ch7gPYGnNz3EVqqypT+BQ08MkeN3DbfAsYp6brx27cAyOCtGHV0o0q/tXqkoMwUMtrYty+C4NB7Q
Y2iQNoFVYcmNFOp7qfFRa1OlpbbED04BNSRX4Z1SP+MN01pLk3UnrLGwXxXs02qTByHm+gE/VnbS
2N7ZsYz3Ky9P3yHWiVjkp25xm/6k6xblJZeum7DdRMnxdELMQ/D9jKk8NdFQwWywb1gpIE6ywHQl
lwFMtC+RMIzkRwEeRD4E4riZBvJdS3m4SIPz6UxAvzO/FmJAS54Db/c5HW/HhmHY8s0N2SHlCYue
9FmHiKy3A2UXov8eRFWdU0xUmBy5JUx2h0r7ptkM4iUkmRM/ySx0Dw2Oh7HxqpnF6LC20fcokn1R
CyGCMty2ZoU9acA5MvUQqCpCfLvcVdC4341QXH+s9a5mLAIIKV9W/4OivqexOotTYiL7aW2Mx0xg
5ImvgmuXzKTc5kVllA2lF9aqV7WodeJydzGnCGZouT/t6NdF1CjT58jc3B5f/jfjK9ITxixYtRno
sbz3x+I3pdLWP4o+IyhS0n0fcfzOOuwwxFfBJO60gnMRJKIyVR6b2DkzziXdjOXclf6TLh/j6xIq
ot4/S8O9GT++qnBGcCCLNwgCHlE6ce3uMNezv5gSKbVWsTAq0d+37usVBhG45fSk/et5fkyWSNoj
4U5IiKAJcLhQsT31ySR40XSsD/U7QJvnLHs+XGJuPO6pCuXwqcR8gdAERCU0ydYbV3/VdXFXs1tc
BEcqHAkr4grxAEf459Y1fkkwwtvBPkMgGd45Nbvu18yZ/j3MlXzbA7kM7zWdrMw5Q6Q2BObwl81w
AZmdb/ovHSmQWcoPan2lVPw+01W6q/a+i29EL2segFBVDkoA4KoDATzeQ68juP/tUS9k+qMh/pDA
QWUq7ruyZ+fE4Q/VmqS0Hkdi3oda4Hs5s5kZY9AqAibFaVuf+FE4/FNkzu3PPCuTKjnwadnPEX1t
Guh8gPF7ya7eIooviFTfKNog220zk021RUUvEnvd2cEwc4fgtRvH6+oD393eFHCWAFsfTiI1KFGR
3cz3xWBKH+5bCg4tC+eURaMnmqLnXwXKQDz/fw1hmtJ/ibySa3Gg8ArDOFyMs0kE9caBPiehQ1hb
oyRARhNveZ0FyzLyYXHhBfocJ4LyDe6VgMOwpFwwsbpCzpoo6usvYdWj6A70CB6JogRgY9g/n/+4
y+iE90EVmXm3c+yQxdqVjgCMbaJtZdw8FNfIpKTK8+7wjte1WJAKAn9VpNsQ42DE9CKV77ucd49u
1v7M+teXJBFrBv8zLWDbBhax8uVbgyMctvvJ2ONpME0NVWbEstq0ZHF6Ha567ASxNB914BSZECdL
i7xFf/uU8hWC33eHIoxjOPJ/4onR5P7qG7dIaAa9FxiYib7f46QyCzHMTpZ4yjufMQIJ78F8Lknw
C6hZ4jw7qZ/z/Oek+gzN4Rs/SCkviulamJEpdPP3AOri84l/z0XAKieckq4TYvKB6B3hkp3w84qE
G6Q7/sbgM5aYUYq1AIPuzZgI6yZF37o02arejQ0eLYalcEOtATIUdDZ6q9q7Qi00WWxq3TDJ+Nxp
/vfhaBlySp19hFFjtpGiWPU5u3BVMRYACE8FNKF/C+IC9yPhit5nIjIjEFjI4eggWuyH2Lm0YBPK
a9IG6//iVE4OtPf/3zq6vLWNJWh00OEgL32uZEXEW1vBdOy+UT9BWwrsxfwbq0nmSCHYaRFZrgps
olleFO/33avu2JrvC/rQYPMnGKC7C6woLIOp7uGWURsgOz1tps+4A3halOB26Y3Zs/4aBG1LCRKl
iMNcTyErDGGkhWa4vA+jx8j2pxftmgBbd++TdzKuYkcjo+wPJZuBFHMgSI+Lkkk4X7uIKBmJ5kfV
KgIgh3JEQGh9MJbENw2FTfL1vmVwFAM5eZ31juoJAAmk24Ot8XamUOt3MCqipc2xPt7SXLV8darw
ow5irJnweLkTG6fGjmLnFcEIVvhztbC5XFenLBJzr034IZNNhhBYPvakvPKhht0zGeSaQJuQ6n5S
OEBzcCs8saDW9Pwpgrb+3dXVJHU5r47FozNlby7gzvTNTo5GucRqdthgTRA5Vta9RM2YGXwy97+A
+HCGNPcb4AP/sUxtdaIMrlBSKCmkhOBAuMgK79zorAhcqcudHfKX06g9rTYdS5NQAFPW/iZI4vZs
GrS0NyfyatgpTfUBtpGIvwYjBMWHpFOd4gXwSANH23mTLER9Jx2Bm7a7e52UBG7FepR6R4At7o0o
kjVo980snF9E3nXb6raVo+77eJXE4XIN/cyoNNve08V4E2jMrrQdBH5YMswa7zgll/GuL0GSjoGr
nqPwjDf7eGHFoQOhpCAhLu5uo3FXBbsHXW2SxdxJFPF/cKLnZe0DqhkLY4DVVlbyNP6YDOa14EGJ
8+Dr9Fgq3WMgBlKVDaETX0EzRToOA2KpuQvmMEyINrs4+symMg8xr9xMB6No/YpL2VesYEf8MQ8q
F0d1RNir4ZPhoE/yBoG/I/HBUCzZUd4fglSF4Di1xoofUy2nzNaU/r2OShCSf18rkhEgBxuYnJm3
fiQXBgXE64hjrD7ZCChvHHRwhxHspfaq43Vmh5aw36lHoUfhehNMr3CVuuXJtX71K7fwOIBm8QD1
iQFuOdHoqQ4aJWG7XwaTFEkYEb47OsenEi0fo7oLcrXw2cs79cNNQ2baNRyw8/oY+Z2kAjeRIzbv
mXEqPTLxlXWmePsUuMetuzTBYctCxIYldSM/IlaRurCLGuj4AWFIkSyjUnk1kbzMJQU8o3BIBtda
phc/7V72h+D8cmovuKoAIE5FXcFK7lt0se2sZex2z6sHBy2xT5wj6LduO50nNobDMNwjH71/uXwh
zdIiRBG8zcSF6uVywVhz7GQLDeesY9EaI3n2vHPxFZ50IgrZMXzeH5vpeoD+kX88Zl/lxLIzxUiu
noae9Co9bjcy/k+Ytm/ne/IYCRJKrHyngnxTZNlxHLivR5YX+RksrZ5g0aVHj+gmQzhHcADE+faV
ciXtQSPvNgvNbmZQ+yJqey7KoHLTR5mhGIilm8cRtHWEyV88bwz8mZj8YtaMTxJvE9JbybZmtylh
SLXDbMvAIj5HiHwPyoxG/q0/ZoqADJtOqbYQVA0TFYesIih3J6Jq5nB/MVsNl0F+RFntv8m+wfWT
tfKjmevzOzwt/Rwg9IerpaDSmGaJSgW7n5UKlC2ALrSA+vaWipEMi+sgpYH7gC6hHOMEzmON29s+
m83aby5jQY9Qu/a7AIqnKNLZFLSAiQB3pLiFnTqdMqarOE4uvSDyCdFVlKYA2PzSjem7+lOe2q1P
9Hepf+xRZ4Mc4qQPQrHkYBA1w0EasScG6qxbGU65JLbPx6MzVPshVuoAqv7dsEYDm7g5s+ZYBAPT
1eVzLNLe00lQ4YnpjpiWqfzduLVudpGbRLcP5oHa535RPWevZgfeqoRPfOkQIo5rh7iK6Ld24s+B
S6bjMmp1U/Q2v4yYBhZjtnaKFMFQQM9l/14rMc6Q9l/49pae6vp1RTnmRiUGn8A0BeDK6FkedHZ3
6HNt/w3Rt4CFN0t7NvaokpTyjbbwxm2HVtWMK0kcH8M2eZO9TaTmz7WWmv3dydxOV+JfayrmozoU
b+ta6vzrqkXK5ihM72qBKMSdfMmncI6G8QZ6UrzIP1nrbH++xsoRaBS0elNotW+nNpvVzLnMn9Mo
cA9zoXpJqSAxZMCfQ261vp9PNugp7RlPXNm7n8hnExQ+dCInO611pdaGR2mEBYA+wPZgjDodiKLL
SOIBSQ4/GKVbAG/AMnW9m5lUnfHoVVUkgYRBoTjHryNoqomp6DEcJDGQYjEUykTYW2HkfKTCLNHz
8GSslwLFrj1adbyhj/L0JcfX1eJjTEAEST+eJ+U5TVXB48CG3iwmSMPm7+0krJqzwCbTxM+xnyVA
pBD4OU7SqJEkb7GbUK57iG/aeqAJz9OrVy72E5bCDmdG4BEIxBt+kXiYcf9QJAkW1az4O7xHbt71
smNYco5O38wDzExi8h/jQ3EmiYLkusXh2QX3My4eYWTOHOIyf1WD7RVxrbg2NWCaM80LpUy52iKW
3t1lE5jT5X9SakJaNYAMZCJG9aQ2zNb8JHoUrRu3LoITue/q/YQwUIpPvF2VsqeZB/QHWRojfLN0
9kd6SZOpfAa0ePgAJDYhr9PmglQqSY+j4uzccxnI5x+v4fkx3I9kZCwCROo46XVzzSrfECqsUNwL
0E2FHsTAwZrJvaY2bWQqZYPdYnhogeerkkPsOOcaG2M8agJeBqcM4iHTEGwYhTOA95UMY9u6ILX1
5YSLqqBJvphWmdxoChah1EtmAXDTuYnrvZLVRk8GWuv/X0mlEjqtVmGJNss1ipHKC+x1coxJTMuC
aswn2rdmTMI8bOHg7we/sLWVwg//QxuduurIfAt07BCzZFVTTbIAQXm4C5QjU6OLYS8xvc32YHmu
Ni/Lwwm5v8vAJXr7nf4eqsPg1w0VL2nDx9YnncHD4vfT3zcbgfKhHjwH3WXN5vuT9AiEW2HmLwyN
iFghj7jgOaYf1+3iNsDsnZb7mgfniQX1OqwYKZsyNzApXTAUN0d4h39N8UiC9f5d7C1iT6XfNBVp
DrcGaESvaF8JMKBZHMLLPiZGEyOVSro1H1BMTayK09H4sy74PqMAJIFbGgA9Y3iOnZt6YG4mmHGf
P/CUM+fIKWCF08iAfNInYrZMIXoFwwZbWFVRIcXgNigdNp2pFrBYGR7CqAJYhGD2czyHPcC7w4er
q5L2jwB6PL/GV/vL3CVXXTMhxlfIAXKYnYC2ksMyhCxPF4NUFRl9tVnSvDmfV6hD2pScTlGokBwq
ZWLYmvmQeYUDSnrojs58mteo2W8z/dnYc0tHjvaV2+0Y3qxZ4jEyCmRwtmi2khhVAoNoKt/NLAdU
69GgEPSj5ZNN13Wa6+JqGU2g5EZDQgq04emvJh8/Sva6UCJq/VM/l6w3uP3fWr4w9AJPPWWr77Q7
O2U9NpzxYouou/6Y0CAdKotC1cZW9NSZ8tdN8Max9S/J59Xd7YXjr2yNJ9s9vGFuCdXaX8LHLIKD
2qdOkFtifwpEDzvmKyAcyMATgKqY60e3wOHsJhMDHs/CJwQNYkAgJsKcGNz7L2LwL7PfK8bW7gGQ
5PjzxbojJFJaWtlEyC+Tvi3IsdmnDesKkWhEiSUXXVzuM8nIM8XA7NlRsd9tDOHLPKLpRnsnd8gP
GA01qWUo+JiwlLy/ULiKGQCrb0k+PGnRScsg78jhv0Qw2La0/Fkma+xwE2PxDNVRHZ4jJvLTR8ge
ozXLkiCx1MUUUjTEscbw7xfIRFpXgZrULvTkmN0y4srWzj1aUgbZSv6p2cJ/rkZY2RgZ+cyo/0aq
qFV44iS5ri00854bxl0Kwou/vDRuZJrwy6/kcWmQYzoxorF9yEqSzPCG435ESR44mUm4Cr3Kjk2r
kgT04cXmOAk9XpWtp7BHyVKY6gApFHgdxhDg6dX4lktOOZNsvLqCVf1VP0Bz+cZlSrxn+IHMvcph
aNGCX2dHQoM6JJ8bxtSkpJg5M4Q6r1BQIAXpYl0Pp1h/4gnsN4XsWZkU9itNBtmovNUJ5HhI4fxw
hhc+C9IqoQoZmkNRE4yNffJJSa/6gp68MNtdPRo1ZGobfNlSyze0szwtwcHpEj411nnAH7JdrBJC
6QsklZjsb4zsNuFMEWTxyLkNMHKniKqEaezhvtmnr7lgSaa5d/QjrGgMmvX0s/TsMIqU58FmhX8Q
vCGbR0ScSrS1wEk6BH3HcAmCjMvloWaeXCS9Zcm72GlHj7unKbCNPHdUK+2rnVjwIe+ppMUiQKEy
3FblW/jYILv023dwOL+Zlx9peagb1yOlGPfL/NeSWx4mBI6VWLxP8VM8BG3QvuHSQ5Lb8sN5pZuF
vG7zCux7BAfGSN5nSdYnZkMBc++YM2upoxKc5rQ9QqHhydWRnaoURBAWMtMBzpvjOCstrwcAeVfV
EZpOh4IwzyeqaPt6VOUvBF74ywI7qJby/xfT1Cf4phZ6kodHr+XbfSNf9mnrl0auzqdaNOJDfklF
hy4lbZ9V8TtxuI57wCurbgz+TOo1l7WODfEodTLIMdRiuVIVDxDg3h+bHkFrIKSX/RfyoK9uiEFt
a9EJyxs3PJalit9CazqfKa2VrUjL7FiEnw7fYM4HFQoSXeZf/X7Tot2l9zq9tqU7mq8MGrRwKu0a
iZg3dKHz+zFdjd533Kc4aLf/64soVVojes89M+5aK0X0IvXYygVUH8aZK83tuqvGr0el8UUUo8Up
3kPuSsnz4+qY5xMTJ3bhNI9B3OlYSpxoPgHg8Aej9epWRC0TEOkhZAr7NRLhsjDZmWuWcb0soyvH
dinWWj9RmW8WbRmIr88RVtMk0codjnnsVFhwkDBa22NIy0M2BCJi0IGL+dZC3/EirBdpdxBCfp7A
2MMS5+bhol8APjeqKdf0dEz0RsDtMP0LxSNg0c149MbgG1I1AH0jmeuUYRbq1HmkyXmLGVpzrWd0
pVSgmmEakVrDjjJ3Aokbl2fNsx6oCyzRfHGOUAwT7MCg8jo0tegOPqpBuj8Qajst+Kzkhx0rt/Mu
fGTVdB4B0gy8mnlbat2ox8e073sYR3MVVcjgeVmiSXydPBmpuRZhCnW++KY86IHgxfaI9xu7HQzL
MABThyWcZxmF61mCz8bYQiMr+PGBZ4gvxlaoxXscBuOZrZpJC/VWQZkNhkFT28uSVI/oooaU7rWb
Ehll1AmWHrp7985iRKWCs23z7RIbAocSeAydSpl4JMKG2P6l1CIURQqt5LnGUYioS1EqFoYdq07K
j7frD6liYD7aXEMiWold3CY0/09bYsUy31B194sNb9qvaWlNxG6zUdqlb8wKptzoa0wwCPtIyiBF
hZCuRa/9SrWO2/xR/FHF7iyXCmNiY3PGUDCHforHtqNryM1Dbl4wsQS7Bntl9SuvNjqimf2nplFM
DcnMD1AWFNcRsjVNw+OIaMtGmxb8B4QVhSVcdYq1aD4nwEOZ1HoDuweiwRvgH5lpi208CRQoKoMw
7TGeZgmUHYqsLkV0jwK/DtwxRCoH3UgfGvWfWdla3D87w2+8hKUUwOnNwxqx2bEuJGcDX40qSOlP
XArDUzTSNcFJc2Apq26tVBnjDuYe5Uh4IsLVfRHluCVVSCU7f3qeiy4id7YUSs6tkce1uMCissab
BkpHfbBV1nvCQ/ePYRPN1/mDK+Mg4gWB0wWkHEznejkXE8tHfFgofLs3YH+YQDQAo48NDO9ENVEj
Yur1ERDnzsjwYtkKRuRmuaHM0e2N51dVSeM6G0NQxlXqrS2rVRV3U6LrqAinOO4so3kcBjSjmNCR
3zhySQuObeVEJPRfd2zeDXM7/LIxpIAYanxodDhIWrK/XnMNsDEmmQvj2gNkw/hqTVWn6nfo5JxC
UeY33ebwTth2Xq7aIdLFvEcJvCxVo8u8v2I7cOHXlDWUUe7emFyVTNTMttVeyVjpZT0TlLvVlu33
1CAhKyv8IpgscXh/X4L9z46eVufKb2+N5Q2hcbrQrTJhFGsDtWZWX55O8Mv/lgcDki8MYgzBXafB
T+CRm5GR4FeRMsQ075k7KKGSsDPlxDpffZ39HfYSwNeQ2QMzW3APIycbKtL/pq529SafwtE0q+7b
Di+HlFYIY6s5utx8CNe3ZkiUZpl6Pzl4BxZxhlZ404a2iesPBDVjmVEHYczRedQ3G3eAdJywjnkE
BcwGoYHxrZBMPb5IwlNc7qZ3nbM6Wgjt5VtYQl3fqIU5n0ZBG5K9liqyXbRwkziUNlsx+GyHcpOz
nerVL91GUlaRMV7yQEfmoFSAPtnfELUJ0OgXgTnh5+Nn6qrzyVnpCN65SkDsU4bmB2+/WRP1SUfe
Kw7rskuSFSdgQSMj0Yu0z+Go4xk81Q9MfH+7lPzQcpuNXFnZYdD765J0t54Mpu3ovKy6XYyd4xTl
vLvzVLhsTaMWfBFWxdDuyZCoLh+ZDX2RTKB0G5LXEbTOQJP54x/Feb89sbb/P3Qocn62mNb12GnY
SwLcxvsnYBaVRldPOTiFC2ZenSUXsRhmEzl3O8bNT6cru+xLLtym+2OazdItoJY4uAjw6KxfoyKk
mNgODm5hrtikE5EPm+PROVj+89IxNTJQyX2mKaj/xWA8/urRM6dmTn4fWYzUVzcBrjlKIPofAPhJ
v5Of/rgCLy5cGH3Q0CYKRMFf5JNBKLhgjKjUCWqwdnnZIAScAtP2V2CRC+vjyjijAlHdUKo0bnQS
e/SczRopBudDTSVanGMEu0SZ70CniJUZKzyaXg6bzIWI151ktbjkQUP8TNIdCX3YOfaHQSAmnh1L
P1FssRUYfhfe5z4I9HX7T5xSvN5IGzI8Mg5hg0gvUGYMvYSmhoxMvdBNtGVb7Hbt8IuOWZhrq50r
84GPARGsz5wtxoK1ODan6w2DKbrRMd0tsUb5oDu4vlSk/cs5ICZ9Z5ma5+gjx8QAc119LWNGOjUm
xA9q60WkDXj9L91QBSnP2tSkVFWR9tMobwUcC4k6iu3Ruh/W6rET8+lDQjHpuZMZnxcmusFEKcua
VuLBKpaExzLNPpkkzyTlLszkaCK5rehelB9az9MULOoeOkpnIv7OWb7gdCixuu8kJDPQXmabPP6b
VmI3JhOp4wbVjAeQ0RgxoMK3oT3yVcW9DNzhJJR29huHzl4KPvwIyDJUX/iI55r9n0z1bg1VYDiq
mCcDBZhT/QvUxJ1ttrAc7AfXkMc7ajPEW2XV1odCvjXlznsGbD7KuMXODnE/uWXoiroHl5zbkrZc
jp4Lq5qmpXZTiIuX8vqn0/V46MYbFvH3qlFC2TwriNvGTHWxALKr6W/QAAHjbDIKOIRpa+4al7PE
yNintq9PPM5cPwuL/0++l6VNM5AZE4zNBdvGpF7mcyU4DU1WdTnVaYZpsqzgF6Wm6YTFk4X+xjqa
Vse3jjVvg9KQoljfNP9buJsQezXVp7+Z4NlIvSkgjb2WJdx1gZD0SLz+MSX2RX5VZ2+N0E3j1TmK
KhdXJp5pM5W9oEtyZntms3P76CRQeoZJ9yzeQso9l3G3oyflat8CwM/1Q0Zt3+Z1RC85yChWJnod
8e3Byj2diSNJCgTSiEwaTGvb9LLFOszMj6jyxhfKK2KFk8WfXM9Ps2GQeCUHJBNqZTWnuHT2ywok
rzRjcszSwbLAc0dtIzewKvwF0FfVT1X9TOlPpeUsiz1TkY5WZ7OQ+PyNkTvRJyluVlNgSr3MR+uD
tGad7GUA+hGq+0aCkjdQ3M1VSFGM1QYE41d1IhCdGgMCxy+IEs+/iFoTXjr63D1O9Rw23wadySEQ
8Nu2sEHl/1bN0GmmmejhQ/BIzgnEqfG/HB0be2cr7wAxaq83YJwEKKwquaRr1UzczgbZLqNXrKTT
lmSU3x6jXAddaxz8yyrEHzDw+uRqHzQgw7cjIoRuzKXTGCUzgyHtdm1SAXJFSdaOYQUVDBeguMjx
05inIeyxLUYXPuc7i3sI/0FHkJSMJPifMRS3QLfA9QRlk26RsTmbWqEFmizq4JR5xMoGRb7CPl4L
CSd/mi+/AeMmw33QTNr/CIExbo1V6E5lVkp9/5dBo4Y5QnC9xhDGUoGMop4h0QrLH7uHVCFDLu74
fK801I3XpyHW2LlzNzenVVXV9SmUrXiL4fns++f4hr6fUPr6bG1KxlFdlORDiGICgMAmLdJp72+u
1ARVzM+B7jJEnWQMfvixKI+52AxWMkWlbMzn+IZgvBK3gjLMyoW3NphwXBo8PaESFntEaEpLak+I
9S6gL1aR2c2iZYkiFDlmtJIzikTGcF3m0UFdw1+MMvaDQizZsDemwwDSTtLJtQ7/X+MPSXK2zjQW
Nl+pNMoLPUapc8uP+lSxKGnsGxehuEhovsgpPbSucpV9dGTvWsTORAHBfEUh5AljOSeutu5vGPH+
4uLeqrE4m4iBqT4NRUKLYZIvjfIPHgbDRU3ek+A7cxZdNyOCXl237WdN7q3K1PAy1d/4JNb8OypZ
/ozmdYmMWfjHIEIqzWDS0HmsQSDn93dR9HQrO/OCkmsaK81uiX7s/Gb4iVT/c7Kury5wejyH3fK8
1x4/vJjUoUVCI8PQ9KuzbBqGhUUBiO35uEVqXc4sg+yh2q5XKzr6wOb+oVqkRsyGAbPZaRq95o0m
C+sXVZN6/zjeffOfbpDhH2taerMSJTOGx4nmyE+2K0i3ZyCs0Azl1YP9RhVDq3/wp77mVKnuaY16
MExc9zEwkSi8DPP6xkT24LnMLSxN+3UfgZtTmT1Ah2zTwzqqYd2D1WJTLpUIEtCTNIF21b7EsBap
iSb2MoXhAmRrai2EJGfvOiHh9QJBrkXD5HD1hCsufVFlxytWIXyf0FuZwQSmkyhQjw8HlwZRxBA+
P9t/fJhnkKqZerXZ3VuEF0ZBOu6FMI6EmqRazXP54LStY5Dp/OJ0ELrINTsWJ3ismhdL8C/iO8IP
vPnkEBC+Zo/xgVSnNgZJSaRDAycV8G7aeF6yofjtTgcgLS4dya+nkv6TX7eyc7cbPZY7ACOLwF30
lDwuW9Nw2MiVPKd323VUx8vI7tWkPzdcIRB9IcP6S/9N4WVBUyfsda9rOi1PcTKGFsUK67sxMh0o
iumfq18SUs6FJulw0hKo70i6tpWESOzzdfYEYAOAxLlsIsas7ByYABvnDyh0Kk0mHRaW1HEYkq3K
51EXYfTbOCbyXNmdTPCoylhN8u2H7h1uLLYPJNpcijcxefR0n7s+fpigXG8skZwRIS63bTQAy0li
qE65fLFAfqfaPXNtMAdfN0VgSDiHj6vjr9oXFi77S/gdxKHYoRuVWhp8BzAH8Ne/R38q+ttrqyCS
r0Xfamc09ko3dIIyqjWYbyDMyFDM6bsITlp+fZ6j3CePBDrJyRM+VluzqtgmMc/x9Ay54JYFNl9u
q4clt3AlU5GSAPLxBVyr3ehAlACUA7Kj4Uf3ymZ7bNWChgxSlJTJlvEprfzPSkbyXF74EjniBRAl
sn5x6PL5NTPIlHpOI8olOkmf688gjzzyPvMvrbDGTGE3pToAVhilmX0DDHIPCekBKjnf56KrsfhI
ohYGPcQg+7ND3p8xhJupFllDa+8RISFnTHtYA57meAkuXuWtb6n7raNrS20DA5RPLyqv0Ftsfrsu
Tb6ZAvTKoes+xPGVuC9NturZ+7bkLkzjqbatf+s1UIKrrWKzrxwdXouPM5SqLHuXlaKHRaSOUIUz
Bc1f9PmDdmYHWm+w/oR2BRg6Ye9Oc53ShoQSTeXPYR9a92GvKpJsO85o5r5Y336ZNcnPRfJAhDdU
rmJcIWDGM/X/BkxACaLsA4HkzFnJ/aqMuRl6iAtUkl0US97LvvMFl0CZyJ2gn9TsUVg4jYGiU/d9
pcHvhezjibKQrljnEhyEX97LJ+p2RZvSdXpJUQtFt9V1aCT5FHKhmn4r1y6hyyqB2cCgyosG7dyJ
VVFPu4hP40ZOo8Jn2lg5igW9LGuHZ4vh/QnbZictMDHvWvU5hqnrrsGF5jGUOr8iHTA58V3NQk3d
3mG4gAsg+/o9wP+welyJ77hyMW0eu5oOPvzADoSTk38kejTOqJRvnSieYc+mrmIgiNjs+gXTUpIY
Hox6oNoLnJxp/8CD9AjgAcXpHGKahstQM0kTr2UTca7W3h+8pkVTKJcbt5KZ6w2r6MMhZJVDfNWb
swIsRfxkPsbkW6YCUT+o81Zstdl9FFLr0+AqeI8fFpv5pP9+QCZbcQCHUnYiB2K1n4sAvKyu2Ble
axk1qkqctn68TaqylwDmjhxnv19QGNTAEUCZFMDYNCiowc29wRtJa6xt6iBD58mT6DlefWSNf9sh
wH5KxWYCYhAfGKORxcQVCy1dzmVWGDeOmYjFOU04MstRJCsLV1pVCA5aKrhP0iiqfL//L4S6pCFt
152yE9E5y+wAT5CvfRMH+zx3VVrzqHnze1RXPIHeWKEgctpdMKY9KnPiEPRO67Zyqg7LQxSZ+4TL
BSbXAFNme5c3lzw5vdxSIwU5cj+7vMxNS4+9VgCt8StnB5gU+s41Sm/E25sE7tzwfRG/Ue2Q9oXb
L6Z+aGDp2jSCg0wu4T3HEtvvRCMM/eBIleHBBbIY9qdWTsIKnBqJxFkAvZBfKcvslECDY18hXtjD
59BTkbUAUzSMMiDMvCvqUUAGxur5N43Kvp3JbsVDwp6LfTdDKTEKKHTK2VJUHRdqaH5HbLeBsUGf
Mb4olaEZIuEIkPLNC5MT2MirMunJ88PEFcFdaR+R7K6XtHVPmGW5D5HdJu1DZs2PvJbt4a3x5ZuT
XZOjSgmUjSiCKfEe9hSbYJ0C+oPTyVwyrs7CHyy0L4GxJTks+HM2r9GsSyNMPfqnezTRWUMMbmFb
pbbmSSp2k1VAh3MuKWNiiDp6BfuYOAVAP35nmC1xSu+5LbuLnS7p0v2SIRaHhGA+5QRSMg3V59GS
Ej0i9F9t4qpnbhi4V6SPiglIvsYUUEaJ78kZ2xPzQzGKh1EXfE5qbTANXD2DpAtAYlJ6ryuraVGO
F5mDHFDYS3Eocp2vHjxR5vFc2/o2GnQ7TkykI9L0qGjMyHzuqYyqwfyANXY9UUEfJbwC1DyLD41Q
cTAXQxH0biqEeroRLYCyFDEXKKb6nys1crJo5K7zBcYG0VsK8njceSY/GnfjEEQD/cS7QhBa0MM5
kOC6N9QUIk4j8+ppjATwgRBs1+3aZMcjWlXAgQGOYUm+ts1OEgegIkS0d5K3qj4Rt6m1IRCeNL7Y
F8UTqOPJV+F9LDQnZapkzGf99EkJhr49jbFmyk0tcIIEjC8L0FIjZIN17+GvVUmQD1tGXnaASIsV
wyup8hSlgj0QOS2xLS+66ryfSJdhR5fX+yWiymuAgVA5P1N/aKdAP+PHMEP+y7IwC4W7aANKuuZa
6zQuwjIQjP3MSPggyBq6MPVlBTUVW7AU3CGPZ8eTHiLYzuvn88FDLnGXe7Q/sfmPIq8v37CbB0rJ
VIafKLirw9JYRjax/2tas2/6l+vTla7zUYHYIhwOSnIEX/fsVwtbtVFEHXJK3+VYWIvEudRanP4D
4CTuU7ebZQW3NyR/Zw9ugo1oCLJ6ImCvY92bR3cEEfSTh2iNVg86wYYXA3jdoVfVp/Ouk3e8F1nd
qeXROox1G9XSNjIwDE5XHga0xEe1wDNnXMHhaSMIXoNsIs3ttFQpvnZ5CTla1w8YHyI83qMsydCQ
OlqxErVc+RJvM47MuKlSRazlAn0PHhpf0onh1wGBN8DyGAMXdHF+8+f+STa8s2jtJty1JH7BuQjF
Crz6GFlIajGv2PEjAUtRcvTiYhTaclj2ZAi+lqtFauirad8dQP4lHPQ8z1RXqZkY3WM9BgULlflm
FJh/rvvhelfXBFJO8odtFLr8sTFxudORaGn5QVVKb//d9ZF3hrzfcPPn0xtS9iQSzA2RxKd5gAvp
2/9Z25TSxkRPSHnAx60TY/gBVq2/ncirKMZKvuQD/lL1d0bHO8rjRUfvBWbC8n5i5L1N4g4Dr3bg
B7gwqPaijo0iCBUsn19I13gdIHLkwmccK9PTpLdI7ULkwJz6BHuRZk16OdG+/yuGnWr12+OvS1lG
vK1NuTIEPcyIme3l+Lg8nwEhjjxDHkyZ4FbsmduG/bSGHdSuzGpipKqr5OCCwWSrnkbq3P9m9KWf
qB193WYOzPsRp+IgqUq2+MAVx6WsfihltYoiIY6m4JGUFtJhZR/GDXsdpzD3Ri6OBvATdHzJNL9d
nnltQbdTmo0mtEpk3NX0k1zLvp9007fF8Rtcu0Uq+3p2c/b+rkp3eZwCARyykFA3UCqB3RHVYDBR
XCfBgrCDn0jaMWnm+/hOIzcq3R/0UL7Fbz6RS7G3HHR/R3A8mR2J9DQRxmSPP7bdqes1RPpx6Z6j
hlBC+FfVDbe+JiNKv9tsmJLzzbNgDsZum8w9Fpw0/XfLaSvtg8A2vkd0Y7zRnMN04mw86xPp+tfj
RPL+BB+l3xHAz+1VcHHA7Nj2ksIrID8uva3KNYfc6E+UCOeI3yAln10lm9UtQ/Ibr6lxSlILkmwK
67t4TIKh+V8KEwBlVvFCnVLXkMWNeaqj7ieAve1KYeJb/kWrrZZfkpCn42O8RjL01X27xXRM5HEt
ORcneOeZ4kbJxvSaB7r0+wSLRlBqKxilAId98nHn5Yysx4RyGXx/xWodVlq0syHpMHIXOB86E6TD
Ifncx1yg+AXzHZEcZTKlNcHXEcOlv0lrka2ABzOXdFiT7PCe3Y0tckMvPIZUfTTfTLwoeNZMSa5n
Wjp8gJHCdkPe6mBmwRZ6GeaRWN1d78paHnubWX9ueLCzWbeFwgbSpd3HzFmspL67uCR25eicDg3S
bf0njdeKQzsKXfHjM+fh0fcBVfV0QrvabLdxuYB2xtWyPsAZZzvv8vbtKFiJP/qfdkiOYSS2A81S
abzyTGdf/9X+g2M7mwytV2S1dsuQOIbfva9TMppIBanUUKa97V2W03eZjG5+tYHj0HoPO/llSuMm
BdH0/4cmUK8na0/id7xpPE4WORnFW4i4QZxzhf040G0U5AISRttGgaJg3K6X+COQvZOA0yFdxcFR
vCGZ0v6IdMwVx75Mm0pxxWDoCpgQ6RxaLJganv+vViwZEAG0Q6v7IZFPcE2bGDuJx3DrEucK8O+S
ewBLMROYDHRyKghi6cxTjlEyAjD9Rz1S1t9MdfAxxoygFgEegVmyCjCOjadNFevshrles+vfQtII
yrVCiui4Pi7UF5/KBK1O5CSvvJ5s0pniOrS6OcN8m233Oz9PmFTlk5VRZfN2gPYP2buUsD/1SbhL
uw12pUIbUaJsJS6us8gzeauC2jekLTJZwxxSd2riACIajqR7coLyljJozlomnnSr6S9V88ikhMn8
ZBZ2exG8jZhW1XZppIoMMAnSMouYsw4XkR7326t8PBmjTfnFnbeFMF3FxpvlaWogIfkP7PsBKD4h
RQ43G2vh3K4qWeepiWo2ngNgoQ7y3ZflFFSFXDlFUgVZSGvsZYv4pXcGfQqsMcF2GP+RAOkITwfn
pzsEBHRpMEBT/Ad9KMlNC0Yoxm6TuQ2zLDq9xQedp5CzqXi4MAaNg7/qKIcSIesJwoBP0xlFq90s
cIvAWjlSDJOHzIT6egwsOj8WrIjnOEpIfMEcoPXR3knGPTRoc6FEt2UP6SfR9de6dWKHjhRYsYT4
v+xAul2LK6aOQzUPDNyPC/HSHk+NqvxNlpz+2FqE6EZiCwR3Y4KHbDFLff8/GLlE2RnHZXjcyPFy
5rtVMDkKVxpBJAF2pZBtbR/0hww9qRnEyY/7J4oSmDTkkff0FPnXlWnsJyyqcyNhtB/HLj2kekBI
XIL0FXX7iFHMj8eiyZA8iVGIGC9CDXDO0x+VYKhi/Ki3AY0UvN33emO9rkGX/nyqzuq0xk+B4GY2
ARG2HWcGIA4j5+acUAj3hsfoLvdAE/VcKuTXgoNMIagaAJgdatA3kdwrOt+fLguiSmPp8XYh9ABk
3yW5jQg0Am7pPPZkdYiEeTq2/V8IF4Wgt29p4w1bhLufqDK/m50cOseDFcKdkkvOXkaKuTteHEmB
7yfI9lE1qykbEao3dXtZ7mwYNmbKai2KzQqF6z5U3067A4WAL4FVcbTyk24TIk5kWVpGBbJKfwaC
feFH4Ul+zSKa3QpNdTIDtXW6i3xWGuwwOhuQDbiWr8vSI1Wuez7oGn2MwVR3B0oz5R6ulrtEVsBE
w+OZrCXzOAvpPuqvkx/uGurnf5yvtglU7zxd45uS1GsHw5HYUPBiP22ZTNGp0NbaWUFtYz+UzTjK
l4s0oVcXZYWcLhGWXEr13B474r78+cug6JwvhwETa45OuiaxXva3KCFLsckNnByqwmMGCVtiWJ9H
IOaBpenh4H+SjIKlHNCrAFDUzJBlN76FrFngc6rI2mp04cu2GzSnkwHCjHTdWhn3Y8NTV9gnaziL
AgIrBNqrGz0OIAFIrplejJmIVgBVwhwOuzA+w7QeqXpIYTzqC3GnKW/tP+AVMWIEUIpBUvDN0zOq
vDSoKu99iGmGouxweS1H10D41GOcD6VPLngqN9pnDNcaHeL5F+OCwNs6U1ZO+m2FXFg6l7vH2HBJ
FMii/4/e601aLUI9FF/ZW1U5pw0ZdhKec1GWAHlXp2ETtc9L+FCaX1w0UYp+Rc6ohokkWaLrOCKv
lRj9Q0jCAPn8TQsJcyivDgEh/wluC2sX3pvIqQ5m/kZ+sYqQb87ldnK5A5v7BCsbDVK6LjFyakbq
x8fG4TPJ8aw7zR10Bt+mOTt0026OtX2fICbi7I/Uyo8RsooZ1cu3Hz96Mqhe0HRJvx/oWK/f6j1U
ABJnVzMGjxzEJ5OU/U0O/dJM89s9iJlEs0sbdtjhXEiov3alD2iATGFT/LmysGHpuc1GBVleS7TV
bqzFm+A20vzEN4OF0zjDn+TF61e698I5SyMsEhFW0/KadbYLFDtPZPmE+cQnwVrdzGHnpa8jhCNw
VxBmEj+veSoi5trH9Xv/fcBThM8kk8z4kSuHhRtmrnCb8VH4LfSCOg0mBcOGeVtK9jiIdX74N1mg
lB6I0EXmTtn51H/0oTD96b4Ox8h29Snk9L0vhmA8YK5jKTxgMCcLGPUdanbJsGsdktekVF3ehdCa
+Q8AY1ifGltVEEhM1bnqczKdZC+yHnRJnzkb9PGntLVS+ObrMVB0PFdDWuOHMHATUWRwdgPfZu//
7c/KJ0wy4gvVP6wIvWcbGZ8d4zbkn0wjHnmWNghQERMwPgpaMiS9zwk2buFtR2nJye/PvuuscMSW
i0WBb/jULOmWd962ytRpZH6cZHQpJX3WkYSHXaRYL5ogGyNp1DWc873Q99p2JmkJvMldIgFmgMop
OL+SHWysFs4adU4aV+2WLgPlQwwDQ5GSrnh3sLdu3QQ3oGdxNz3D71qP0N9bXklOO5irFvnHnFnr
pEmPBdpU9EvR5I/JWdFLyQpCfLe7q8tkamZ7V74lNfR33/qXKNtF5JLFir0Bzp/pFcz1MR99SohU
K/9Cg1+uzf49IHose6VZWgAI9swLDRMBdMYqOX4agwdK0QJLksP1NSbNIAlZzM6qQeIdhQ6EHQU4
AqDFLvR0xo6ZgnSx/qELRR402g4xixgczwxKUW3fEv8Wb+Nm15UiLCm06MjAx7tDcwzigsDosyAj
HFdgkvkiuFkl2xn0013Qlggr8UysQf1btRY4097Vouok1TQdcItrg80jFiX7YEiM5Zo1IfR31ozm
Mpw5O8zXAPGWBIgtdLG3OZD/JRdnIm9pRfZjVQkrSzM9DjisdM4raClZ2a/3td/nQ4sdF0C2PduG
t0uKmZGXhBTgKIzmPWYzFSuRBaMBRDCSfNtkfEJUdVKqipn2nyfI4w7kMF9Hol7L42fXL/uLE6QH
rczWNfTIGvL5pqcC0bzyG0ok+/5ReHYE4KDTLSxelGwZYeMl/9M3rvpq5/YI95YNsCmbW3jLUIkN
DHj3+rdvqGEOumi3zzJma1di4SJsd2sf1gNm9PKUROx2PJv5KV/TJ7C4kpD0QzZxSQZgrsjDQ6hr
ACmk7ccrtC/LKhPRKRTi7j//Af4xBQKHf3kWWgMhTAUYcNMPhwT/NfVIYZGEwWIZvlA6yK3MXOHb
w3WT3rWxKxNMSBM4oGb/wTojIwb6K+VqEoYoSUDDn78wWqvQ8qMz/RoyjduQJkdpnZzJWowPNCng
ljZiLk3dYkHGVfA/sjaUtmGpuD9W+fctnlXiSScZNPA3NKuIK/E7Y6UI4SSN5dpb17zhIRyut4+x
w59sZ2QKBNyOOPLKpXxqjI7O1DIYBZ7TLDOpZvVLxJK36KBC2HheVs9Ui5I7qTQoxkE05Vf1vbPa
VjADNciFKZ4fTjrX8R9zCEFZWB1dUkbjzbQH0ycJE/jmKwqiAr/gE5fFTCsv4Km0eGLZ19G7X4T/
WO1miO6fA6QDLS4wB6jck51/BHfRUCN10HVAOqG3NxRT24bzI+30nOduHgH5l2KghlCPl/why/YV
KVsnwxY+/0xoBLEGlPMndpsqPIXXVH+b7ZvtbdRnRyHz6x1DI9QNeSr1S6SwLAow8I/4sMCZh3Hk
gm5j7yy+kgPPCEBHm9lz8dwQovdHUYQb8Fzm6+hC+hEbuNGRLfsmY+QwQ+nQ6cjrn7yxAnvF2TAY
8erT8bRZnBxxrKFWl5bPZIlJC78BFa/APMCksYp1hwwQopyvTofYyXqunyQXDurvooQDb8pbtCqc
g07dCQ/IoTvMfHTlpBJA969P71P6CYYyMHdLgBXyjgK+qqI/Ps6fAZC9MESVIJ819TsLDDEUuzaE
jrd4oUALFGifrnX9CGu3oQrPnCmS23AHAe9qY9LU9f+Fhi3pJrms14EYzBdrMgi1vWuDklXTYc4h
Z5yhE7uMy/g2nguDooH2RdKymy7D2bCODFnLifm86TpY7BcEiQAkmXDRruazGsSFiOT6Qk3cxWqH
nyrHKa56psboWuITRj8in7vrAcsdi50z+5KBRdnQi5t/8M47UrlU4fL4EaIXaiOJVBdmG3Hi/wYP
VAi9HEUa4GpTe0/2kGQ2mOCJ5wgkaq5VKat8udbHRcwQ6ld2WPgzvd9eZSYsNquZz29QMupUtQnO
7hC5m6XHDAqB2i5c9fR3UyPatHEdlG9CUJ2p59B2J6mIv5KOjPEV0pvSE+kPRmZZPjIVJOKHAQNy
B+5YfK/4o9/W14DNZunQZ/iwRN0rr4fCrA96NAc3w5hUMyNhGDB3KFXZt8hFFoRdHOCVsUOPc9PA
l2fgBjlZ733xbYCh/8h7KTL2wCorU4mtbeuKb1385WgYGG+BKRvMKEw90bE2K/+fchvGbqRsi3Aw
zIIA/mpblq8FCtjDETZ3kQMQFHuymF12fmPvgK++baEzYfMrMpYt7xbzoyDwvWDP7YJdlQQvuF6k
RxfnvJv+skIj1e8PxXryLu377W0KNFkI6NO0PVn/K+28bl7g9vHiunBwnBoUecF/vGoUmrB68IQI
ZHOspZ3JuT+BhWP4ty9VRMNnRI0dEEQNYZQ/Vb2QGhOeFug4WTeAoUYnFtzkPx1VBwXGxQT4MJSe
3aihc2fat/DQPSzfSFYVF9So6NK3ZVqafwtAOdkzLYjJqLTbEbAOa69MKgeKeUFzZSeLBIT71PE7
avgxi6PXPBNIHEOdmWzVX5TVm7EaBScLvPSOaVvNPf7ehiZd5t4sj8ICI94OIqrChdvsish8zjOV
rFw7+lniSy2N8j+RdZxwMs40+lxYRrC7NWT7gEC/rm03+tdo5NZWkZK7Uf78vGjiey4YPjt6olcc
aSi4IS9/+e3BKE1MP6NtLonziLHbHHmr8CzB0vAWeLUStdu0fheQPjSLsAG4x/xfk85WMIuNI2Eq
iCB9XdxUvxR9ocR89+FwMez2uDpKmotK7JbWXgTB07fYLiW3Z9rNvgc8/exIiLJhk/pOsKKc3HGn
qZqE+NDNCo9YXiyLdAM7sbAnPILUJLIUwRt5lgftxWdmArfOSzVn+KM35G+KddY+Wei8EOwSbAYf
T4O4CwThkcc2P/x9G8w7nmiI4W4cKQF/3+uqyprs6c/YJUviRa8xrhDaK/dy9JWtXn/HQKSP0Jdi
WZjlJZTbR4niXS3XZ7J7OWTpH6+hNmKHs39YxyzS8v/l3NjkDN9tRjJekfthWk4ZVX6C+m5kfXFQ
ZSaTW6X2EkGpr1cxfCJHyDsYEWqd1ANPBW4DR83nkDpT3s0HKall3ohqO1ClMYddCJVyeLB/q5Im
TmSkw0dTTnm8USy0uQL79XFeyAiYxpmO1Uq9HPAia9b4kkq9D2/r4gBeCGs7kX0tmdGS1YQTMolh
16HPD/jHZHjVcBbNOe5kfY89GNF3NuxlKXC9h1KHurGurJAoVBMeCeGYXlIx8qSYfU1b25U6Fx3A
TeEUpXbynaUSilGPfuSijGToB8SabuXUfzU/SZZS/Jy4HwECwSpdFEodCcRWx0W52XkCFlwVjTHG
0ZytdOJjYJ82xNb6kkH4VyYTxantbomW4638d/LISQK7wPRXyvZ1qECLFeo9iszEhzjMzgD3X///
CXOfBJlL9wIGvGJBx+bllP2iN+LxNo45GDnQRcNiB002/Xt0CD91c1Sg/pQt3s8GPENDGbpz0EEz
whTVcrvbdEfnK4wP/7aMqsAEdykGHO2As8wY3w+VsvD4PPi/i0T17JpCXsitHNDXTGaxrn+q49en
mpZPwIX4EFz7U3QY5hUD/9Fj6g9UCzgZLmwb9A1QK+unPNcQJzFMrMtyvj+fax1NNfnyE8TZV8xN
vw7M+uqzrSj8syfgH/qSl4b7G8IVNmV0jrxPjzrG7dPkY3im7OvlwyuYSxLwRiFAwy1QU+XAZBsX
1dF+AWdMaDMREccljNXLszAJVrgEl9rzXtes46YOyu58Qq6SJmsRuWX2lklxhBl/Zd6ned0gMe9j
RNFxA0guR3UOiIN0ks908rcuLRYtgeYS/o+UbKAJ9mhQC85bH2GWCGcaBCIrA4zDy8/9ndnI2TQe
tiWLwerZvpWmaWRTxdrRnPMHeOwjWcDejys3I9FpqAXeequo66+p/W9p1U6zoi+wCpMkOQHS+H4u
0XZHBurIXMwJXef9HjpA4bRW0yFtM9qnMNsTa9CA5OEJAtlYCflO54fcdC9JF57PM/KPn+FUshNO
gj+CkVfUnIq3gfBqpLckbl0CYaslMx6JmMs0pBI100sf2hciA9w4xhYDM/Ix3YVUkziDRSstiwB9
BQslhprWh1nqMN2nRPP3qds1aHxVi+S5dAsp93xuj2GvBy6eezh4ulSghkkyeClb6wdizfOgUaZk
Yh7fq94Kpm0j0kc2D9u0WfyVhH/g5hJ82b3XVpJWpA1r/l3+ngeNtRwFHGJHJg35zxj6Jz6mkjXC
XEtGMVpU4xqrIS4zcA04vgnKCSyN9EPsku1dKWidvkTv06UqquvTQSihxhNgPZTZ3s1q0YzqU7c8
g62PE2reZP0t8jJM491zSidcOuMfiZ/A3yUE/hXkVM9zoExDhuMhrvNsgX8Jpt+bmBFs1c8K1Myi
XchsjG+qGalHZDWyI2K5sliQYiZbaB20iX9t/swZgX7JC5CYm5Ziu4KdXY/yctWhfZm1zMdio0y9
hix58TKFoDNxN4ohDp2lfRMshboMJz0NQ1dXrfqSglAb4AnQLtZsi+ujRQMT9qV2rfaltlNDaF1M
Q39n7Z1KQlmmwq+TMvQRJ+HFUd4LR31P6WRIgInESzX8ORWJ3ux67SWKz5U+22fOrh4lyzZol4xc
peSMmv0qqPoqrJy1NJoa+y7unYf7AoAWGkVOZG/fJdQ83e3IzZx6tc8mLCljAQLvlaGrm0BUp2YO
zwsGEQLWv0nrJHJ2C8opUmdEClnx1UABsoK3p1L5OdceWEBAHPrKAA7NFVMZHxiC+rlyWkhxWVAy
4HWKaa1JsH05trQF7kHPP3mEMpsEOqlXGfcNoYuPaDBOr/W2DEI27seNewwXU2pVtGGVRp8PhbIC
m8btIzP7V0LG+UdK3mS8UBG2Ftco1gA76SfX7or82HHzvP/VbbuleZiqXmL3Qkm7731oPKHhXPDm
726kdQ9co1/67Uuc60XfT+mvuclCkCwEvxMksTHaCSCuBrxzbolh1q+VIv+cvZAfD5KTpu6wH8Sg
ce5oWx5udq9LJ58YNnV1rm7r0v3VFtMEqVJa/mAxgIUICNlwAlJZj9DRvfrRtWUSMrdm+lTTPAfE
lVV7L2A5ZI8fiMm0L0CL/tNASekrjK0BKInCf7NZtM9SjZjSY3yuIlDC3VsE2Q+emoPYvOj4BPU8
pqzs3ElMsBOIYq8SpWu8uAWYVcyipzPqsP2TpQibGWfcFEKnGCTMLc0QI8lvu0fP5wcyPQDw7ZXt
zAW1N2rD00QBlTaoE5eyChvzt2EkEIRodIPN8U04DH+yoe5okPfqxrjJk9OoQSgF043NSzsSje0f
N4oplZvZFuHU7ApjMb0qZnwmKxpd8p8dweS3rXblEGwVqaDOV+FVQLblcT+HvNNkGekm7tW/SPOZ
FFycGPjRfQyViuHZI1wSNWdUaxKW2ZbCdw2Rm2ANlILg57yRq/20tXxKtWDNNS1fGLas3Bdb+IkP
nIMhZvtf7tsE3Wn2mplf5mXhxuVH/AU9ZdHFuSrS7Y44+t/IsxZQ0Ag5nYyjsiwoaKMtjCdfFB+D
KWMrbAVpFDaEqMDlJF9t1Thb+x0eyo59uv8677tqszSArT3PTyram8H7PbH46P4dzORUOODOyzAa
J8C4XqJvxKsi5S992ud3mw5MRi9c/ETd9nw/nwI2gaAo8J9SKm22sw5FnT3UhUZnWifuEtQttGXt
JATLY64EAPPvTu7+0tAi7PKK5pqzoG8mIEMmMfQwZ7JTvfL8BRWiUQVfFqJlhWjf0sWZjrpa6IqO
Mta8vZ1CqKtGKkgq+NldLuz2iDRWoFac9sqYinkNgXeuSJWDK1pvv+wIrD0ASpTGGARwjzKFhh3a
ae+ZOX8Aac4n8QWF6BMvcz96W5NAPeE9l5gB/p7MY4YUKqQ/OB361eg9RkWFUvuzK4a0bOQ2gE/p
RjzqhrNZ/syxbGLlVd5lWGXyXdbO6qHg9Q+z+qPS9hMeHAoxYdlbFHb77CXiasoJQEwfsVGeGBzz
6hKOH1etWKyYmyuf0ziogRVjDvrudBj9rDJYjmyqp3/5IsSkq+msLAr0SeOERZEiYRLbT4tDv4ww
qx9ecUzPf0pK2/8n8vsJHqr21qWSWvgEnq8tK+6TVZGc0yZYueU0K4VnKpMfpQ3t8YFFyDmy3GZ/
2+mGkV3iGH0gf7Z8OJQwwg8EGkY9og/6AVk7bwB0A19LUBO+Wzv4rnV2hARZaD+C5yMJN+IT2C5Q
tpmYiUXFp9qvvlhyaEbYrr89P6qT4TgP5Ib++n9VykX0Z2YvqvZQV/X5BLzjUeZ0mnfDqPfwAxMY
H/yguCStqRrWt3dZRYVikNwl0b0ZbWQXymfYSsU9XmZFQuy6FpAeF8AALpfFzUmpN+AzkGKJIA8O
tJ44AOypjOb1rkJdpBXHUZ7agfb58Bw7Rz/E51JqScH3tJVCZdOYUbf3m2WWlHBZOUk+zscvNCA1
FnjwhQGfIJIsDFFERHeMjoiAsUNof1rRcUv4/ECV4eK2qhAaJBNcsKI9dXHYNyIQXoo7K08vgcB9
jprO6Wla8XZJ63jFLF7lWGObyALsCBxBFjoG1zxWC3a9ZVJV10wq2qgbTz/1pRwGH1Abj7Df958Z
h0Ur33JjrpQ8rnXOkLBzFFIAi6OFkkqCt+AwIk+mvFCtrDQxrYxV6EQMUgLKM5PvXNbsoN4pphLT
jGW8vH/YRsgxCMnBsgGmQo2nnansElWaP5MKZCmFmq9U54JYCKJ5mAAU6/b4zzi1WPtbULAzMvJl
NMF1v92IBj1YC+RAUzPoy8/g2yHew54xuMPq8Fsl3jM6HAGahgZn28/konGXu5DkPdKwQyqWIrwG
jIGzaDD5QdVjOBcCSl0jhWfBGjjWWFGsFumjaG4JO35ePLiwuXCrsYy5IguIPZSqUhU34H41Frtp
pXfEOqTG36E29vYjAWCVFDid/adPtm2vB0LbStvD2G+zezq69XA1j3hOUMYy+LNFRdZvh0h570zE
MOKnALAZyo5yhj5EwdBkWxOGQrzyglQ8bZ+4vjwIkAIhrVbTR9H1NPve6sDN30BdFlUwFBIR3BIe
xhxWHZqVT7aK9kQgB1gakrglCZYRib2HPD6pDkBvg3hqa/RMArZYiWIWqfUONiGKbp7KQsY+yOLo
xX6A50m3waMOTz2UZOUIBvIWvuCmKtjYJXt6hgNIlwGKx4J6FxHobjL+v8HW3mv4oyHLLOMedKkB
TyFv2wbPBPAVTLuYbRU15i9BKccTo2GoxyWN1say5AfoFBiBpdj6h3iFkuOp/V6EJvfd4S7XCNYh
aOJv18eavMdGqX+uMW8DdBkKFF0UXIbgYkDbzqFT5t6kRLe9u5A1NXk3eMSZYlWrwAEJbNiDEujm
69RGpIzEffJuwl3XNTIE3Nrw0QkblHQt/KyM1PebZmGrhRTaV2vLCqNPQ85w9IKbSem2RnhT+NDa
ZZLcCn6c/Ncfynv5BLq5i9/HXIsicGrj0diuOs7FhQaLmk9RO7JGFSfxd3hicNW3K0r1qoGPixwD
tUyGNCfjOoLbNFZqbnEoFZDiW6TiFJXMtnwzwLkA4AIuYFw2H8Ke/5rBVwEr1711HfJnkKUXg+qw
/xgB5W+D9g0rBa6kaWgzbrZx7nsTa8F9stQE7L/UVXoBHRFvlLgCUVXKXJhMO3bNbTTGJQ0QnPLZ
sULikEdTr7TF0xQW7q9cGkygn73CMruHH8PSJWpSWCGs7FCn5jal1ZH83ZUPoPOCm4uZkokLtI+I
KHh2Gh9B1gU4c+A7grj/b3wTDrXQNRLRStVwLDksxwTKF3z+s9GXlR1i0LrJJgiRlbRSICP3P7br
5ql46T7xXXUACcWZtaoSXph5RsDXDEa5z30DdcB83yytbg0THE/H7xSFBQ2QnSkSIrMMkd8s+Rqa
bKS9ww+qYcLKWI1hgMGiY4CYwOZxFzjPKUX38jNrAc+48xV1gFxZl6e9cl5ZniaJr045h6tMkT+T
C3dK/vhIoY5bdrZjcLyfz9rePBUps2TP6tIeIjrno7A9mGzgz0Yh98fTxCBdCXsPYdXUGIUUvJmc
g7nMOZNjxxpbdCdd1dkk+roGkP635bb0FMijzx6LUOGugp0j/sODvcuL067kuSbsOS12Z/XO9x3U
ZmE0cbEl0IeF9TX8DCy1junirY4fT+5x4DSnCKILOd6GF/oCySgVCe8K84YD+cOliHwouVgh1Vyg
YCxHRstXzfCtYE7Y3OA9AXjSk4VH5s/aiaSPU92QsYxU4b77x6ORhEoM5Q4XEoLnnO1bdjGfpDGE
Mc7sRL9kACcGIJ/BoM+lvrSz39LiMhDm7Xw7sYUdzVRsY+Hz0kUim8goYKlOiwdsgTSFMWTWqZ0C
7tYmaLqkqMb4wgVqCo8e5nd5cpfL3yqiWDE2BahAgzBoRhQKpA1oVJLIOrOd5frFotjKk7hNXgWp
GxkT7awJaZ+aanaHSLmBwmP6npjUE17mRHv8Cvmwv2Wlpwhnkl+t1odcTTSlZ+3apYGdIP/Gljox
yPcuLdEFj+4ARS5jEKViQNPu2EoPHNlSTrqG2UoMx5g5EBeKNOne7Wb4FivSCbBwK6+aYuH4zhoT
F1ZnTvaP/QslPP5B+WgVD5zKcmRXKMGtL40D/PBcYXElTf3K3hC9oglvDnMQkiG2R2yvVXLXLqMX
B7R7BXWI0NRrHgu3/bUJO8w+iSjqSXzSQYbx62/MTQMveBIgXZvEcK4Ggu//AM/8clpyVGNO07W1
FZduqnqSTwmWs6coz+fpIg/CvwUMoJsVuOp1HG+QXAv3wR5eSHcATHEu6geWiKCL2i/b05jcEagF
Iq/6msmH99NvaKpzphK4rq29V6h71dGRU1uAcIpGE7RmXmdwrPOLUFkvEuDYYxu0JSGepPdSUGRv
Sa9tDBSlU3GDED+/HKmkLyaTtybfmm7EKZnegJEf832mV8lI2H1pGoQBrFa9jo9o8cTfvVLQ4n23
/G0BOlGWpO6wjG6EeTZ6GZCKkL+s2R2CjyWCA7ORYYEQRX2LIeE0BoBEcyIG6aUTW0MFuV71VI0B
/b2TmURhm2HAmA7/YicPfoYM3ZlE7f/RKTvbcSzX+GO4zbszsFPlfg33+2tUBuhi2hNHCjYjqE6Z
PBK1+ztSLpNWVq7AJQ5/rtPm0Ic9sdZgRSoOrtCCkxUEMxz9GwgGNV98dB+RLvngAmsNmCv8Lkqd
iVnRUfIjd5rpAz8mTLxtNDL1HvMKGzbqnrFVcnFXfUrtudoUZwwC5efzJ+OihMPcErO7vnlaZwLC
7teZaU88zG00jciOuvvbCTXsSggc3olS69kMViOPUvTI/b9/zpO/CfobFKXmW8C7flTPIeDo9vlU
VmxkaCl9BtexCEZj16DNO+VVQJDW/HX44kGBug/vXLYWcbSM8JlzqksMa2xs7IkOgoeBDVWkqMXn
GjdPfAZAMHJrPe1jSkma3N0V8+4c6/tM3n3MkVi25NzrY3t/51ipqwEOQAoshlNgxYyWAaCE1+bv
CUHK3xbgi+wZ1UDaGKgVRSEaZyxCeBP2QZReQmISmOsgN9QMyhvo+uR7iJyetMMqHgz4CwB0rHUF
RJEUxfa1jY+9j61hf3CvQrTIooMkqpXngmpwiWGSdXZHTXpIb8/hAgaS2ONMp1OKWjeyMUygmbzZ
b+TXUUZn9grHTeRuC2sVF+qCsY6pDvHxLcQZUV75QEw8DuPOmT9eQjhCFu+4A+qK8zqUQ9XCgG4x
EKrWsl5tFww98Ebr6uTWg4PQ69/+92wLYNyo2wb42HWK6S6vFPOQfeYKFvdOhDkJl1e0vbnKEqX2
w8jgMSjR8p+1ZQqZKp00N5Psed5cTIkt48AQaygvHBjc/rXzuPenfB1qi/OfCMpofGcxbNH3NTK7
XC0z7DrSORnnsYItqqZfxtdMvFsqFlUwGbKvRTXwlRlFLOzeeQu9Egxx3f2+5coFWVITeo1vRcFq
bKfwfT9aiRBoCgOl9vlqDEUJX+9vCdaPtFgPsoyLIV/4gtV2ItLVFdqGUZXoCMDht+u49Z59tc/u
UqVUAiU8XV6XJlOdZnEBIyAh3nJjiYJyHq7+uuTU4sB01ympQgi14O3LjLC+26rGoxBgbCSgqwsH
U+/R2U7KFZqzALVVa1ogiNvbIAg1eZZXYUof/Hovq6AvSacKV5WTUabQegrqPbi/LWiA5BT+RVnl
QoNMPj5ApoCt7PqB6rGkzyVJFuzBbR6NWM+9ymeFNTqEZfUKPIy4pQGwEQC+7vQKgDUgLEco3nSb
QLa/AGqqqmfFmHzL8V56j6L0ImMkOCVIGvq3S+t0phTWQchxG/lCBVRd9Vx3fsEOmL/OJMMbWiz9
kD3t/Po2KTQTEQSqMh989G1qdA88zKlMXTl4bqUoQLB96bSqWoNUE2HvMcz23RmekoZMBcW0KlZv
0tLlxeS66GHdP5hJRwOCU4WYjGmEp+oiPGVb0tp2n9aaRjAmtzZAvbnRRJo/vIO5VFONUP9Wx+P7
pNOKLKsr68DKjf7HUUM3PDOl6RteZDaN0NHmLmaz/3WQqjvXYtXsHY2weqaK3eOGgrtnmfa//cYR
KAt+gxycXCL4/inYIHBOBMiy7aIp25mAC8TRmBkUeOrkaEb2eSRZWc4mGZyCZrxMRDBieNYWiSmT
QqPehSF0rF0Z+VJeDflAs7/iPUQxMjJK2UsdQfvbcPpaeLDwP3EiKol+VcWgZp2CPl/8oVOLTvm7
NN8ZLVSq3jBftk3vwafUL4tnoWugeEFIOqzsfUo8FtfrHP5kLltuY/fGzrFn0eenBfvvgvPZ8g5g
VL+aQncPfrVkM4U9gEZqmaDUSPSkw8LTiy4cAd6wqJHhSizYuU8Dwqe6gpUYvmTIfDK5WD3uzgwh
SWYSyEkpW2JNwm+N51Uodx9UV3ftkPaoqzYUXLLLH3wqrvVwVXRay3f/SpIJj6TRNOZvlSzyTQty
igs0wOLv5YHrVg6Zemv1d/6cn7r9NIwM2t/74+uuX57IqSsls2kB/dxLqt4wegIQz7VD7DYpBrOm
g0c2qWL2A21D/HgfaGtQPP9/JkdDtynV6m8ioCs2+C6apCMCmvw10hkT06hLKxDy3KX6Cno6fS2g
8ac7JGijYqCvpfEPJmsAdyIqlKJmclC8AcLVh9EzzJy37Q+H/ONFrC8QAtBR6rRcmcQzeTOA7NMF
zMrgbwSM2YMogkBDadEND65VtB9xLtRBQJBeZU3lUuC/7sc/As0VxmqsvbhXp1qfyVAxWmxxzKGl
pJQZq5IALqkVtnc4nR63Kbh9G7uzsSnha7sB/cm7TQoUWn+YSwjRaU4rRggmmH6dZYpfI9s3CGOY
cGOPtwJTOuLsbCWcMaoNtoz3tFsEqEimTtIpznBTEin9D2NlZcU9/sGBsncDo9GV7rOygV2gRzdV
qfupGqv4Vqe2zPracMt1Be8XbifdnvDjxg2IAG2tSBuqQIESngIInI8ggLFVw/P7yD+TQ+m6YLDJ
zMwiVLZUxMwlkDfD/oU9Xy+3qIHxxBuhLUFIAERIGg5MjRC74wkM7CdZsULpjPIwYAZUO+YbipLP
aUxc0+iW/5K3Yxkeyy3MUpUwxfqxpLVMN5ih3WhJhl9/WnqowsOxEpOjI9zwkd/Z5Qhyau0k8vYP
nzjyl2Wujjuyp2l8ZS5SPQf1jOnhoV39uWWcagC56+2dVoyRqfboLWN5j4yB4tfHopYTT6so+O1p
UHXIzvwDjPYvH+kMXbYOPey1BSHc+lcmIBhl+xFv/lHtQcFwZ9EKbSZHDkWmbrIk22y80QeQC4Bb
8JLQr0CBjYivZmbsIhSaXPaEMGXlhy8BYwG4YX5syeJLLTd1ksuRr5rgnii+JTLi1+dHbH1qz8U9
hzblKzLnwDZ0O1tF9TcmgfxAI0yVBLsAnu55zn3SBCrzyWRrLOWJ4ysJuBcInEYo/dR/LN8s+NGL
ehhgYVO6UjXvq+x3ovBjLNHPFSgy0iDGCTqEcondEl1yYdn0+DPV9V49juAsXykDD3vnCGmZ5hak
9xAZ8Jhr5id58psf5LVuUuFeGFP0sEzVBbrR2AKqJC3UldNk3YcLAR6xB8pxnHev4vQD5RUGtgRT
dFTUHcployN13BBHY43ea6vTY/XhDeSgRTFGnedVhBQxHrwcQYcWQKfkHBAl2wLIoHUV+3aWRB8B
wyabqTDAc2vqQLulWgXmMaDBJMQQKHSANbdnsQrLSbpJNCCu93U78DoCfWuaFfdrlSDa890EJTCr
Wmipiu3TsQxB1D2pITvsR8tOFLWwDKSuaTiewev+cJOruEyiOrSmrTq+uZYcgnib2G30+GDejhyX
Fo5Cd7JPvszFaSq4RaxBD8HvkDEX52cCIImDIVyFpqxwAOIiHYdSxr/eHVt446z9iTKiAOCwbLqU
fpOPIQl1tzYHqDDEltjKlrFcXklDchIAnHZQ1TH6MH2UeDZtfTf1WEOnDFa1QYXEp9wgWwDJXGHN
WRRVdf29kAyOlH8oll8qngfngYQEQMqjXZ2+m+rkh4ehu9wyOSoFfL5A3lxZM9wmTkZN3uVz3wHt
3N5oi25aEOeq2AguG5O5nMbxvHfTRLrC+KiCUWp10UHtTe8hkteYvRCumaupWHOf/Y03i1MGZpa6
94Fb7GJzaf6LYDw36ZzEqOgnfF1ESjFSSywN4IL/Cn8dGp+lGivwX9oNfqWyYkt7Q+/JW9TTh/68
Y3453iDBXnr7ktAMy3aanyLE3CCctQX3PO1DGhXI202GxdCdOYXBrVEahcOFRvUDQyOzUiYOXakf
w6TaEc3bjOOuCnhcemSGQxnCagxcbR+iG5HPJ8xT+gdxN4WqAAi8S8+UClFPEbPkwHojOpNigVVn
CJTX9dqlJ1KzD0k3agPjchcAZljg4CHTzMFpzPtiMiKYROkXMq46FTvnd3R2Joz0p4zCnXv3fEIo
vy+wAKWKXCzZOMX6JzWR+HR9ysyvmTyUWBVY4vtIGf7tMKJUPxfaDIuZXzqyTXVD9fLMPjD2BCnV
WQd3rn4Yl8CG3oW/FvcFqIobWbH6qZd1ojDww2EohnNoLE5vazWp6HbPy54413wAyDZmPgAD2nR+
SocRpJYt0oELHQVAgeJIazppzPNdQaGeeBdV6dNfndJfrZLwHowiH8lz2SprXacQP6eRW1+gmmEh
hkA+a/qhrWOUP1sD90o/x5zVQSQu8CY+u49rQlik5d5fctMOPJZY1VII3OcSueLMPWhJkGDqrE+f
hDygWZ8tDINOZABIdiac7iLpKd+GRyHf2lQvaOoCK9F/qeDI5IjdZnLrGvabKOUCFa4MGMKlnk60
JsRyyKvR+Yd/Sdrhd7dov5qIobEkKsxvJOtkM5P3FOu+F9R53hjiKDATYQvwtkRWXnhil1x2ZbB7
c/YXdcE+hM9VwJJ1VRkqCZGa1zbgAlGQ07RFqPRn7LcD6OIH1s8LpQGwoZMekepCsanqcajImYUk
7S3MA3J66pTLk5NMS70qP8gkDh+WGkj749kpzjYKtPtFKvqtWmzTg6DUrLc6rjdm1OUPRSyhmmpY
LP32ACWxd3ausTUQyAZYZMmwBtDNZZLgykrTp1p85L8Fcp0pO2kwXDIEdFcvDffVibq/y4GIzn3Y
9l3V5ilNCGuNYhyJDxiQYSPCYlHvMuRWsnTzEHZALuaWglRIq1vjYOSR8dvuBDZ3+XEA8/QvdZgQ
W7U282Jpg+5nW4gew564aVuxpjl8DbyMOvxAmdUu1+oTO4HqHCpZyIxKepmJz1U1tstrxBHjn6YJ
gQF49RnzkHrORUY+lg/ZdKShxwXSwGGRLDdcj7zByrXPIcX6FDTy8euC8aa6R8rUY6tSP591rYgJ
ePQurJuGHVxZkJCFdubVoUXspoLgsFX3bWSTcadtvlIXwHbiBunNqn8UCb+MtlTLW48UaIn2YDOd
br+XZ1HHQVMDAsyOfAsa9SZsVAXKKssjy8rn+PhhlTCt6iJDjHQChvpyDzwmrXZzFuPjVdsfNCE0
2xxHGIS5ZfXCJYWEQLebsYBbC5YXavenMfMgwnVvEXgn8TxGK+mLBwvPM56aWS8xMQpcPXRNI9HY
oyDjb0iBKahE6vW1YqNVF3dZ3CQaX5S382H6G672nHjRezSmp0uzAT6eI0+/F0E1ZCKiLINZzhWg
CGqdifs8GKKvRUPKs8EqHX7XNpNF9W8WIrRW4LAnFr2knZXU1GvrQN7gXnwKa337WaD9ds4p92+f
4G8fLcw3ey86WO/ZXusvvK9PiCNp0Co4I95DIhfnc4nw+ck8Z702SZHfIG5dwIBxbiBHJhCD5HML
Nrgx9OmVAejFSmCyfks5tiBAw6zlvb3SAwLHPqjEFsBdQ5knYpe3RzH81aUtN5jESkj6ob8M+hpv
8PHvjn0vaB3yTecTdmnOPowJrlt6LLTVVUp2fy4UkcrafFqEFDwNyELV2XqNLr+gTGTweQSf58zv
grrTbL5jMDVLD6kQQ9OFxZLdJftv30TaC5LZEsqgCn8JeOeLVffOMb+rbdMkaFyYt6hKbc6Cx2kl
6k0zNCEotWiLDcG4ezom9rf77xPaccMG83Khp5NPqLDqXCR2ooUvaWHNCdAzhLxQWqolL9b6rv69
u2/cz6YgaXrayrkySzK8p7SP5hqQqkUjxeXhWi6JJqKiQcEQ7M6pC7T5EClLeHvFEbbf3+k/VsBP
7PW+HRyEseGn/YmUINZkzFoMFy4oFBwHg3uVrFXfQcB/UkIvn2FeiBhTJlmbOmqItG2GcZGjuf8F
HYs8DXHdULWSe01d7EQUNZWBOPkofhJCxuzoy9BTC4YA6Ql3lOFm9ubg8sOjWebnfN812SMYZohw
psdMz1dq+POhlz8o/dYkZsp8vBzQg1EPuqtdAq8dQ5qrF8uBNW7AGDiK7BpyZvumSbWyKF3VdBYL
ytqYrQkVK/hlbvoZfdbYjWE6Rxd9MnwayQIo97d/ajkJhJsOAC49g/9iGCo43lWpET8rBmBdBd6D
qcodWuPenScc9OjbMGDK2Mp7+ZmuuZPKejTTgyM7y4+pyTEtXUy1h1/v90j3NRBqiT7gFW7AW7bT
ipgVNdSmuWpKnc+Ueh0M+iBeG70lp/rDCXYIOkncQe9Z8MyHd4YFOscJ34AuHHiwqtOA1+NQOBvw
+b/jTBH3pQaWSjAYiCMRJKD9QntPLQggHve6MOQdhUpogOKN7J4bJRxsygJnKVMa+J+eQyI8AvDB
7a9a2ysKFZzHZvRlpX3AIqxUNyPhgVYYP3u4+C++0iEZVVwS69thwdsnj9ztVEAwru9jgp9f4jRQ
PULHP6MhMtmZkoAWcbQCWmXVZDvY7GGHT9I+DIeiDoVDygo5VctE0925V2/29RTATlYqiagvShac
HJ0RtEAn1zFxFUXffsG0M8pb4qCiNuQGhbjXQfeo492Pl6dVP5F3yUE83nj9DawDRw/M4GQZnqRT
mNf0skC6kfRqW7DeoiTRN/4WkYlZTJXAcaFAeLBFF0RccaTNa8NWcu3kGGuFXdqMqvxUdDZCStZm
5aaZgn7k5uJ8lv737yf76p6sRqxNS2QwBV2u/XEbCPdksKAjC93l8U4PTjFZAi6ee70DKgr3GSmz
bR1VkDNUwg87UNBDkT+Co428qVRmINlo/XySkUcFHuqzIO47K+saavtyo3coXISPfXMapEnJ/Ldm
vqobB9uT5Ghd/ijoPAblvqTxxjPTQ6XWLXQ0E+UaUVrN6lgTqifDbsik+uCbKgxrmTByscrMc8Ra
ZYRW4cvwZJdZcbHUtf6OaKoS6VGnx3BDF4YNag2LglpprQL6FSwBueKuH/pR5Srhh+FgTb9PWzPw
vxtB+BYEf4XO5U62cXzII4q6vZltOByOGbG47KI3p4SBuhLi7q6WeOxMV+uDEPbXCnf+72oyoZ+Y
5jcngXmXLhkMrtd+JpuHudtSUx3j40pe3ZMNiBBrwZccU0K1sibGuYr5+3BaS+ZQAN9EcEn0W5qm
fCLWojfDwGDZAY6mRflHMo2IqHxT6iVgdargE/tKRZd7/zuQd51ODxkVg2OPzliiWLGYdftUMEFM
1K14f8TXQ6oUzEnDJfjWdaNRuze5EyKbnDbEYqk2mtcZQsCYHQMKFN6NgZR1cCzPdZjMb8lne2FD
EopuHAXOd3HvxAwvsdaKdumZ1JQnQH/WXO4bz7AIW2x4c3SOfePhXAcyKorX5s869xBiq3gAJmmi
8UbS01tZcqwxBNoLcbv0xzRHr8OvRBCzM19eAW9WsIWTpkhAn+RJjGLmwyzdnO0kH6ANEAPW+Grv
GQYIziYNQ91n5VAGbac4KAQC7pl2N+4TofnObXP4GKn1SReOiwTH7Xl7gbjkvA0WVgobwNgHYjf4
q+jRp4+hG7d0ZPoQee6xgjqSIRVPc1MZ9wg7U4ZxG5fdIwCB/us5bHrn7jA8vMQdkX/J/lC/2s2N
4fkL3f4NApS7gHrd1e1a6BHhrkk+oGfhm73FJ9jZf43dlAQJbzpCUR32ldzLav4JgqVymy7zgNYN
/NAhOLEqKPDibeeEWRczSLAO4CVflOBM3z6andjZsodk2FgstBco0VAG7H40IW4ZtADJ8kVAbiac
yBEybA0ZydcNL90Mu+8hvhrvnFQQuSIVJLrbjCUFN4CoEu17Df7bfPPVQ6dCmRWtWOgZN7c/aPpU
E0kDaAWorK+zL6X+Kq9L9cxZj8mE7EcRiEUw1zBCkV4EFpV9vzubCMMVdi8CZc+ap+FA1o5Unp5D
Qrr1VYDRkoChG8QRoimqm+yArhwZlg34p7txFq5K0a5Dphm7IqdCadSOtqvY09/nWVRo8833AFCV
rtFt1ZtAtsr5eMadFip8zctCfc521SA53eXibyHyNlooxE7+Nxu1gvm27xx4kuKRlQA2s5fqalir
QkvxgarhkdLkPpnj/n60LsXCU+zFPAMpOCGdV6DhaeKpyem81eX7YD1dglu3LJa2Ioa2Rqd1iKGb
y4yKcTUuETS7tT83WqGjs31Q3R3JSwqRa3/K81r6Yqmhg8+bK/rAh7W2zn76l+2NN7WF+EkYK0ho
mWlHYnsvMxvmTXxVr6FZwFvnS7+tP22wSNZuR+f4Zd5wDw+D4QVqdPYo2bW/H9ao+ACdse1rIENj
aAqnC8KqQ3AtLLcjIe3uNlxbwCfAP+r5U/YA13KAsmUwQ8K2Kaj2jS1oug5TQ3CojE9D6FqORhu2
/xjvOIRLhfZ2kSJgCNqjqITzpgGjxnPzeOBEQIqlK+0uqG9IkHWcZ20egxmQGX++5lxnH5vdlvmu
L/ioFjgvghSy2UXUzP+490t++mlxtdDVv9LhHWpZMwK2cpw8I3G+hh6P4maqTtvpJzEAlCY87jjl
W3TctUgTkyGy8G89YyPfrra5/Q0buiygb89vWiDVfiTemDAAvzNPERrN1ZC2y9udlGeoFgf4Qs/b
mgcdqPXTTlVbAnvj4RFvr19TNlmZnlWgixDxeLcykft/IFNaQTtXu5KvqHnwXU4DBrIIq/T60CQA
JmEHWdsGCyC6VcGRneTJY6jwUhHMPNloXVOdyAnybjX/7mMXxURT69Cnig7rOP3cP7LlHfU7aDJ/
K3cJiETXeO3lBfpfZZhRS8bjzCYDefSpBqWnNLYqgbE0iccY53c1EcqbN/fUszscvLFtatx2GWR8
kEInRtPjj/E2GWgfVQLfTxMTmJxoHRG6V8+VBFomQPwgHthzojITBXzrT3QOyl8B4u3/OGjnzfas
akws8O9dkt0GcRoNVGjq4+0YytwQkkx08hwFpE/FrWh8l2KUHaiCpwlOOQcDjdmV3OO0Y05ymICu
lSke2laSLnCRtw73NEyWadLbWAk9vQrUOpfryyxZSqCJy00DET0o/pTqWt5bN5uUI+XdGxp/4hYh
tNtfnSj5n1hYzXTHNBctS3FmOBNttBJ4UpU8t0WTPRKTEpKMaLyoW+yggaF39HEkitF8r7RKeM+Z
cIH/jWiB5ff472DbV659FLxNqSCwPabP4o1IwZoXe6A9ZueqdEIEbDdG+z0q4Qvtmc/fUPk4j3t+
G9xabvDaO2bgvQ99fZzgfOUBgneK+71CGKBwx13LfEDNj0Xr23D/oOj1+hpG3tbQq3IvwvKPJxd+
FQnnVuYeBoqSM5lY7NQtW+WNYJQpQkbXVreSf0O2XgfL0uo1FS1z0XcOTAjBsqufjug5sWl85MzT
c33udqDzl7U2S31XV7sWSADLk+Ci0PbXqVxR/yEm4YGs6qwsyQSFQHkow/jIrOFUNUwRQ6KrP6la
T0vcBaq4dp0zXMouBDC3D7GuQzZFbvDTBnnlVBEM2HpDKkiqkjmL5IIK+IWKjvf+E9RaYFVNVm5U
zz6TU1V9Rmqtdocs5QRl6esnl0RJs7RLoe89wvreEU9xFZsD93nA/Iz25v5d5tvtSc3ZC/FMvTrn
UB0upoNVFT/7puadT3si4gTnxm4dCwQwnjevalq2pxyhKOZKAQC5XSIOrD4KAiP3IvF60sBWIE7C
80p1wOr64KA18ou68b6oghWDUbDX87Zpnlz+ujyuvVExtA6NkHsRxkn5CUVfv2lihbPr0xvAFs4f
xLaLgwPCuHjQczbk36KUhsqS+dEMmI7HiB3TyS2lj5WfdHTDSmpow1UCCtwIsIfiUnMHc/NHTX0A
LGvrnXdHF8vFDz2/jnSnAQDsoZ4AttEqUTAnXdF1etJAROq3kkbiIWypcpYO1DfehVnaufzgPq+T
J7O/NIwDEo/oj12aFNVud+jfXji1tMGS81ycI5ouWDWftKXoQitAWgRMY4X13yeTmScozznWJWEI
fC32JNoqEWPcDAqpoOvZRUEn5eOhjeWYShyHeXdnu1HHQql6zXgo6mHqDJhILgs3vnlsROxM0eOS
fPsZR6qHbogFEBKupc23q2dZw+iTo7idl3KI2iwldc6OMiJ+yLpEoIAvWEB3FrQ6XeTQmLhzHARF
wy4dehHzUUlVQCkP8K3KaIT9sbEW9giNAwUvIwOCjyeM55wM9Q6WOvWddJznFC/nNRUQBBf2bwiZ
85pl5Ql7E8jeNKxqXAb/XvXtM72nIK1NTSd7mq7JpVXYcJW0hehoWdWucxl01LIMtxTXcyePdSH+
DH0v0CSQd1dc9Be9v8khcu7eVFNKBE69wSxG/k1Jwy3gQRfPYgac3yjP4QToQT0rj3n6t9LGPmc7
0koo2qPE/cJeuBD/Aamn50L4Fx2LyTneAdIfM0c2ynHMBlradgc7Oz8nxxUUUGFF9zg+RPMqkVBA
k32YwXzx+kVhidKxuMGzYuqI2BVwpryHjt049H9WKI4/8x6AjZAt3tsRcOb91oMO2Ozl+vyvSmV9
hvaRezCb1H1nxQsj2yqR3st0NXyhG7AMWY9S/ThEfY0xCYPaSydGr8CCH1TRJQWTOBIxTY/xAzD7
YLNkKNoq1qr5y+4ACwDBT3coWW9RCxOOyDTOwmHMffiEVk1UyJxBgjIF/6B+Nsj3pt4JgtkR2tPH
QIdp+V+gupC5daXhMGC5naldKikBDE9aowiMX+mIcpmqYFx+D7yBWRqofGVRNEAocufexD5q1ove
IATXp8oPh5BG3qY3ebD+eVF7vf1MU7yTKVqRvHx+bVw7q4L5HiI/DDWIhnBSeJo2I9GPx0V9QpGv
O6hJgkUBKaOfjBRB/y2RJIWHt2ucfBvT3B1OFuM6WBHrlbw887xObx4iDNbpMlMW8AV5kreolGM6
ma1MgtLwn3JTFi9yxpso8qDaDMvWNPD0jytRNrhwwzS4mvyWSxpcsXsc7r6+DchvS+mUwD8by2Wk
cUPiZwRMp2VLQd4BfH3FH5ZTcjJyGlrZDDbtp/rH7r/j/KeGGG3U9ihTJf+2E5VYhEbTo5orewif
WE00ODgSLgb+MgGuJlIuVlIM8/PDLUq4e5vXcLXpjJY17Olpto3mT0qjKgD5ev82KJCpSB6tG++0
Ebn1AZN9ZOy/IIiYBRvqsicClHxKGgH7N9E6PGO6HFzCPBb92WE9Dqxmnm822e+WFVJT8FYCtOke
XXnkVH+9tnjEGa977Rk8CAxaAef2+2+xbC2Yxn5Jwfbtho2xbBDe/+KcRHBkwczSgjOgFGMz6puN
dT5uqpvwNhZtKRS71+PYZQJIKxDl/Z/xWzE1hraWhwmFbYmvqLPnDnH/eSP6fxgvfx8rR4QMaT84
ex354bi9FSasiKDC48DUzDdn3A3BJ+YDzgdBuOozfiL/tFm+k8PwS6/VDFKKNBwka1xFNZAkrGrq
mOlpc+vt6QSIQx9MtZLNKdd7p0dulYUb2Df1vxToBiWNW4V9PCt10uf/vaRI/bTMoTmWJjExytwF
S3W6z/AILp9pFrAFdfQWB7lxrgSeN9tFLGKjPo8uoBr0DFdAXOUHaQIe9dT8cC3BrrUsMCUuyO3W
hToMifru2cEMKVYd4R4Jciot6GXz955vQRqk+dLxvhVq1Zc2QIldqua21v1D0XVT6qN31bEeOzfR
LMXY5Z8jTEnGXKmY1gqh/DIkijASyPf6HXwXE9j2a5B4MRvaA8PwcaBXon6lx6FmDFDhx3eS2Wga
JtFwHn2jS+JNE4xwVUI+5MnXB+/QFw2/QDM3zEwkQ+edFKxA4BnigUnYq/BmBFwKYxU9CoqKyx8H
HOqv5jOB6jxA2Wqrf8kKozYx2sYvveyFedtZQfCOWkGbZ8D95BBfGfjHYY1KTNqTCDnw/Z9/Hbqb
8+iEZtSyaAVWFeAi0Lz+oXjKRRSf3faTNJQH3vaJiZVD8RMLi+9po+XXe44r77snAmuuRPn2j/eL
giFciKL7rUzvuG1wzlow7BH5LaPfrPuwu75u7EQRKka4HvB35zaoeiWdUSd3Wc47BTUXGMgvqK0z
QAsP20MYuabM6deZPDq5t6DwwEsVZsqQ/WZiPG+DWAvenVJc31ZSe250EbrQQNyoN56x6BnqU07i
oh3yK2iWqFrWjI+mkbFkwib99nzAGpA/JTWgGimGonVg0e0gLVNEYNXsVLvECxVVv0cSSuk2+XGg
MIMbRG+9XIvqAfLS5agjVc72lrvzjhVsOacQkYuP/KaUdeFqzgq13W4dGaHMwXcrkJcuXLidZFHA
tI1v+6RCDi4bnh6q1tyoIihPATyJh4ppO02RciClgf5R8o0JTnE/c3WhS3JqKjxbmWPQqhvGkRxx
sgZJAB/cBquhzgPS3w7XZxqWKSCkCs9Gr0buRVVMKTl8YxqabsNcWo9YA7PXC/3s0iOdojmLxOku
yzoD9TM+OdTXNAwFS35rL+Zt6YOr9fOYQMdFue1zPTzXvrf+9D1fgGSAcRnivhnywkngGldgbPrW
igYF8SYG+QFaut4NJ0d4C/rwt6XBvjy3ZCFAaUz9/ydk9gaiX/GQHVNAk3o9AKInzC2gjxHu0wSC
Nn8rMPDvbnWKOFrzhbwazLaz948DErTlHqtunn2Ushm+VtduhxlmWrNun5HM2Dk85SLuSPkFmWaT
XClGdSMsEsgapxDWk4FInm5kJXH5p6Ql0xIZwc7stRKmx8pIzlvXGKASieo64gtWgIqk8c+1efYE
NaBI4AXChP56IbgXTfAYvB+8hdalVRs1b/jRhO8Lfen0CsGaesG6yUyEVqUYUI69KVyJItsbBb28
K0nGFjXsd8D/uvO/ZHxoS/X+2YJR55UXo8hagdVZUpXDXPIbrFb632mjXuYpa2ZhB+zOvmHlgcO2
h1LM6I2P8gSJEL1zRIhC93gCX4S+CM1Y9mIf0cFq2d5d5ZpGnrblTpLiQGCN2eIOta+Dy3/42P3X
pPCXIFGJ439znVwbJbSbrt4g5BOCTVrqUfP5Qr7K0yCzSAx4sxcY6PGmuZ/y5l0vK2+cAz+ewoLd
IJLnjSNn7qVhiWF2R73O6qxCuaZZURDV55RDsbo7WPEHCYYM3vZCMCDYABS+/hHLtuWM2QQ0PaEa
n+c1274Ez3qMzUXjggqB7FGyUV5fdPH92FdJJr40wza2ueszh7gYmP/DYF2y6ktmAgiFcFqp55KT
jqTx9sYDuu866Xe8GOa12wGIVV6oU6v350IJMdxB28DLPA0I3nyOCaJgTCqROFstf1wC/rzSyygt
ISr2HICjMBZ2JcGh3eyNtt1K/hulOJXS/qnDW0G8/5f7PdQySQzPR9uHoPni61hRffLrKSSo2Q2O
hZNvsO04rdM82CeYTGpH1M/ytXmk0WIkn5ic4Qd/QP0sW1qKu8f30mVkuCrT6gfOuRXkpL/Xfbjk
x0uprIR+WWkIsTP+RtbPiyQl5pXCq7so4C1a7AAtMeeBR8RqlC0eqiTeo0XCm6ZlGsLa/yiW60Q5
2fjczzEOUDVU+NaGJpb3fvn75I/7UTNC1s+6PT4QHHbp1zocqsOXa3M5n3I2h5eOsb31iV+CdnPg
gOsywcgi34cs8edvurMhEmQQsDBpRKaHXLph6tlOGu8B4HO9PylHR4SnrTpFxNfHHGCQAw9q3wOm
CueT7t6Mz6NfVhsv4c1xt1DUse4KcdyA+PwEzs+VZOuTRZCjuZeOQYLulZ8/oiSgNW1RQyrqi6x6
GdT/OewzGuaDZUZO1RWGBMSlXvXkFPmBN840ecNNn/q11ruZiZrF2xyEkbOom7xvTrHCSE9bSo+K
gbP/OnrHCs1il3N4BrP4fKfoPQFOhApwGtj20SMvFekWsj30tuziycOdrZgbcfBEMymDMe/6z2q/
4X15P4N0Se2ID2K0p7/CTI/QC+bvSuyclwWCCD9hWRSdDQUzAVB4RgKsiGIP0ra/fnKnzRS1G9CR
UL9Gx7pl/kSTOwB8omX0MeWS5dcdW0PZZftWLp2qathwMmi2q/W/KuWQRxeFbmWzMeJxvONuKvCe
/258HHyKM+7M5OdUP/4TA9l90PeKsvc3jk7due/ckroj9VFinDdEgSNMkYBYDmLcvRnLTUtVC+G/
eCZsO+43lRtXiGJswoscmKb1Q4TA/eBXxuDXWKY0TbbKzjmTg3Yx195M8V5w4RkAjxxk0Dfl9HM8
jR2U3YIEidKOULnuJ7EvygahaEva1A3by6yKtR6VOzho6obViAyb1ergzmtRy6/vB5X9g4QG6Sny
g9fY6gMMZVd+CHP+K9HmwTugBpfrkApl4btAznaAlhJyiVhwErEwHfFddoI8F5qEhzUb9MqGyKHj
fH+jYVtmJvsnSLdDFUC7Yi9gzBBLFII8i1ISvOiTimg/redQby7bJEwEDpUUlxbQxud7BXRKCtwR
x/u70ygPsNOoPRjG9A2SX3AMnMnfDgJV/Y9L5DSZ0ldETlmOSr/Si5ed/6CbBUQTwp+BZYhH9Vle
rPEDWtKuiHwa8jgB+MSrtVsvu2LLVd6bO0jt+3vti8R9CFpd46dx4CLuTil9HD+wgzKW3uwEBzKQ
4I6s7R5A2d68xCPcU5zQPJDKTsH/y1U1yY8GT5PmdtECXtgRfQ61iqQqm5SeZbEjbWPaWvWtjRLH
a/KCG/b4UDCf9ku3bUwNC00if2msTblizmZ0QNQCYihi7ZJUEisGAPU3VrpC4Sk2jeP1Gpf2sQxT
atl0N93Us/H7uEreQxPbU2VkdmtvFU5jzXR+beqpaiOufIR5nhdEj47e0A/ts854Uoy+bH8jRfpa
2fRdHdl7z7q/O4RcRVwDaRogCtvn6o97Oh4iDttLAWD8SnuPRgVYSE2fOPc9i2TtH/ZI0dil5Qn3
3JNletvRwkXY/OtHBGKLbmnITBuB5So6bP1KytXq0BVJBJTsFvegM5r4Nafv4KfsYVgJiYfjehx/
/rEY6x009WkVmVajAx7zw9e3ZAF8H22YDW1vvocvfgl4KyifTlE9dsHaTYObRCB5Bx+Go/r0sOyF
CLbnUjTbW5iCB/wJXK4sGgGf0fg61NNI+5IyOgkWBhIFiCrg3CylT7U+H/XXIBSDrof1woPjIaqA
gojvLT700M+HmWHL+fVM5oeF7Vms0BG4VaWevv7Ko6uD+QPLgXZOxWMUzY0Y9tyWHJfnHWFze6lv
AGFqoDr8ud/5pfX1VmQ2ZMl8Apy0L2ewWEhgq+S05do4k1R4UGG4mwiC3nBO/n/IXWVwJLhb+ohR
bmkc2/AJPLP3GJa45AAyNUw7PRUInC5An7LTtDF2uCjsjgtAdBDivVlLZrh3QhrPwufohrPOkKxQ
MyALbeY0mIUWC8HRpNyAAYqebSqwLF8DBiUhbO4v01NUm5IQaFrI3ACAQAXp1Ws2lMJguEoopG7t
irJzSU1iohpaC/jx8HUPI8dKr5Gv7p24AGSXOfiGYNwU1U7ugvfQBZqwCzEOeXn0f6m1ZEdhLkgS
LcRD1bHIxGmD7g9FZTA+NkJZxg72eVbpC3c5FFad6Wzu9ypDdx95ehT6ohZa9NU9zbHZskR66+lA
t0wKBsB5ClV8GtP4ES8mGUhu/n9xzURvUPn7v+nsphXLD2E+g+9l/ylJikuHkKRPG3Huhdi/7Dxu
wn12pkQhXbhXXvtP6/8cASXB56KmzmU/LxgkIPqXGMOxX1GJHi5o5q1j6Y67P4/NiwxmL3FsNtso
xIu+8Tt6gYuTg5VQYZA2HM3sYpLQow49qOsKrtLdS4QruSjWsYstkejZyOVxtsek9J3pN1vR2nJ8
ldLT+vrV/oPHPpDNzETbtVwlJbqbkQAljmOrO/DrkDFIGUEyT+h1c9Pw+tsD/yzmKLuMC58KG8iI
aqKv3OoTjGk/1DFLF+GXsTKY5ojRudt7HVLuOJ0HYY2eRNGFJU9hiuG741dWDsMTMRgTTPko4nMj
MglXFSGILA2bHzYMqObRd86r4FLeoM55I+5mJGsq3bkog9JmU3qXi7B2xNP1+Vj51Jy3z+Ha5eJP
QFCJxyLdJvJjSI2P46Cvf38aCC0Tl3PDcPqbT9croxSCyzz6P+Z90FYiNjCpI/dJBVwjhGF/sSOa
jcpq+Ay09tALP5iIwgN9DOyruVPYT6yaFSfOxl9kAm5AF3xXZg1M6r+IMotRFZifYAP4WvKwoFcF
hER5cyeQU1o1ko5TE2/SMyVyl9pvKc0+AoJtPrekeOnAiwSdqOWTJzSv6XTOEjiw2xmVVIX4OjDU
aWn9ecxaMqOH0bdol2+UomDnYWewc4vM8UUSKMjTiVCmEPY/uW20uk41DFdiTl84ocVZUeBcwrVw
p1v/5ua1z2r8xp/iYhQWn+BHHs7+a8SqHqSY5DnsLKwXVONQXgP1+/VBW5MRfGDROH1fpEn06pgi
rktUWFdE18NZ8pKo6ELjYmK3oVKAI0NV2UKrgjEO4CfHYaSNCZsA2FnOAxPH4gxmzcwOszq1SmQO
ulEpVxBjqCSRS/lbyCOVnJF0rs9RnQKbEdB0ruoMU2TL+Yw9PNGzyQwOJwkw47qR1vnc/weUVXcR
xqxIALW1XC9wB5SOdSwJ2TW0IytKBG015tL2VbcgGvrDZe/34cKpruj1+EnRcFGyG3FKV+WgK5nA
qzVFwy4sCWs1u0Wwaz7ifVKR0W9Fmogi7J4bqGT0wu7DHI9K1O9yCy44p9j8sJYkczNMCcQaQK8F
2VFb6WlDGziWIQ/mIGuKlTbVOJz+Axwn4Q9oSj4i27ZQF6dwoQmOzHOCaqjpfgu6x3STJxSQo/+m
CUXwbXeygoGWP26q3cpOD0pEfZxQLNa/HRm5L7iExCjmcnBGos2NZm1ltstxqmAivxFB51ISrr+y
oAL+GCPYfqxr5Jp2FMXsJDMcsgNVQ34gqjRzHylj1pTxZ03WifjBXGVbobpSXV/HZA5e4U4UPmbO
rAENDQEqUby8vWdBp+xcNsNJWIzU90Qnmmu1ZVIdabJrV6vnruSb9SEulgeFvjWm3hgQlpDKgojU
UD7fC60BsUrXOGUx6QXaSra6I6k/6yORzyXIs+0l4w2s4ITPfQTyRIn/ZjQXjKAJ+3Ap+OG4S4nl
CZCxpEMGz+xIYld0AnU3X13uwjroqlWI2YzP3tqZqLHQaEQFKdlQ3GVBsFtpzcFOatgU7JvpTW3f
z6ZqAR2bgpGrGfhDBhIJboMBdYW1ATSSvFzCRmZNL4araEW5FMA+35uprs2EKwyQFvVLwcVpns7s
L/zl5BoOOVY0OAXLS+OOBUgm5Cn7klFb6EtccLF65huH1H7EHrqjhOEEwMugarmX18jjtyhkw68W
jknSO58U/ErDxxyE6w90Bghw8sq9YLNFdjT+iJq5qGTCRrmNwv3jF31g6p7aYSuqLE5E8yIw74pM
np3BoE9J18/nMMoYBcZbkVTDYeDiF1IPmuGsMiDLQA81a3a7Z30kIkIX5OWOYgb97RlT6IfqmbXZ
0ijXdQg04kky5jgNowNtRiNwgm+1+fG55s7VEpbFz3DjR2g3sz+MXaj17nFWIpd9O3iresIrHiav
MlSr/HqGMA/fvKj7CsTymADQGSpHlaFcYgOaoa/u89Ia+LLgiT5DASyIuPHhz+Xm5tzJ8yw7iBlz
ustSA2d9OrntpUvVgUsMYAHtrg9oZai+473s7JYEpPJNTli6LzmvFw5UES/eA4nc2yiECQX9lQGH
4HU6cRa4s2J5nrXwF9LMwJ8ibNOf++YaGw+0PQiGuFkLtKh7hOJbGJxU+sJL5SKNm3Dy/JWwzwJX
j4iPxJJ7nVYa/vCuwy1TjREaA82Vyi6Ypc0gpPePQoA7oxo7kd7If9ALtj9jMHYmxUd/YT0nWqMo
uCYSKJY7OGoK5DzQiCnzjUY4XLgazINZLzOvQqNp0ZG65GyXTk1CrmgNRRLPpPSAb9Mm7bcw0O55
eHTpZ63mt2tg0JckMAhXd9ZBKgVXVGdnmQJixVrqPkdoV0cUVK+3w2q8IxsKcJfBpZd6ihUinuG7
RG4COlxOtGOQ66KsJ0/ZqrQ6vspAyMraZlDL9CRpJcbD3sEcJOnyO2+VyGBcvWgL9e7+fVXEZXBf
+bETlNJlskjOb23uk2r7WQImtp/kJEWZIQh9QTaQxmAgTrRk3gGd7UekswJGW6boE4WwcuAgIbGd
3x8fhj9VjHr13jsnsA5fMSlaMaqrNFW+66+k/SaQYjrZwVHEuVQP5It3tH4GnRuBvX6ykQliPfU2
6O9EMmV8d2dBmJE9lGL0Raw5GlREVw7dfLG7Vk8liw2NVc63ssORiskjbsXCokP9VehnUdaKcg/i
L8ZIbPRjuxK7c6EFDZ0gcPUTVHVLl934uNDhrg1oX584PruKL3HvFoUYD7IqRpKE/3gN1ej3oon/
E+WfWBbFAAbB98aprkYmttAvFO6CPp86Rn8lhYpI4Xj0MzPMZSdsDvYqO26yNxHr6NDUTy9k+ggq
A7ySAO9eTFDhbAzoBIfNxY+ELsq6/4nsczMb0JTEppEBwlwOStLKD8LC8B82t+AXZfqaiFQyznfV
RDNXyKs0T4ES62GUs1d5PhZ4I51P/HFXFznJ62c6YhVOXzAFmRb3M87/gE344tvuXQGXHl5wHqOM
Yo+nhOdjqGCkbQKF7RtX90r2He11SUvAB/xOpKzI5szBZ5/Q7Gfy/jiOG45pnXHwyGG2rJN+fjZK
9vk4JrJrCSkjnhv/stOrcxTyv25JETvNwDDPaOUQ39UDSpxmhzwByg4yzjMq9h9gmD5mwwsXoRGP
UGzfGouj+xD2KufiPBeBHQGNTUurA3GUK/jMjSscgZKL0B5Je17Y54IZwJ4Qcr2vNIACERmTgRor
/JiAe8XFmMzl4U4sT7iFnmxFGDz/IWVn0wzSdMTmgz6iafQqhKlXQSjbaz5O9LFsLtI2DyFetD4q
8+fX6qhIr6Ju1t1WKRcEBH2mkobx1PTNGF5wef3O/rpDAQT8CCqF1R0O7bPomoQVXMSrC2W/mi/I
Q8kv3xZRgDk0pMQQDU/9UUo8fyR1JdBQAu6ECZ25qeyD1PwoX4WbfqaT1WQn3Vwb0IHEj0PeusFt
eWafCleKaAH3ipa8SUtx9JRtWYuiofH6wMm3lE5zcq4aALWNx/+I85vHFdPBpP8tmSEVPNZ9Y4u7
XIPEQMlaSNA9skibTirZ7U2pOGl2zaNRXlMPsaF9c+UAmTWka+B2e4HMbt6s3GwvlF/nscCni2p8
JmBsLoDzMgaQaprpDCQMPrragWe4FFZSq/pUtuFQuHRn8Z10J0Capkir0yT9plTjUzND9BSRPf07
4l0nlyaLxuc3EEtn8t7BPf+SpeV/eOzo7C4DbflkA33+6rVXwBybu7PZ36xSoi1Fhf3nWWZ6+STk
rbVgPgtHDw4/821hDji22hVljf5wdUC/BSHfzmQYDGD43Vcyb0y8oAuP4UFCA5XSgAxSgHXlS/4U
hJcbvnPmYKt1G4pm2EESI1YlUFLZ4+0tL8ZBrKKxZVinzvr3ctRevpSkhiV6MJomO6xb/9CmTQlM
9C7eQXW6nvjq3SkXnY1og2xgRkYg8Yedz3DnNiTv/STAxd2tOaJMoDEYoNDSv/04p+y80nUnwE4r
7jpnqUrqokBE4IYDEe1tPOhmIj3V3LuUnL+giu5+kZ8jjok/xbnW78ivEf57swOSJsNSmcDogV2g
Bd6w/T+ZY0ITUr4MD49BRGDnZ/UCA4jXt0p/0k5WSTy45XdVK3d3755IK3kIN7VCPJHymRY+ttj8
oz9RK2q2Leg1rlgJsC/yHqamXufkqvYVz84UKbsLjynFNUGQ002jXugT2l25npumz3Tty0B7z4TZ
4RdyYUkSGmyACR5CMuTSEZZ/ycb3u2/oqTmH3g5S06DpqOCwNBoDlqHIaOGAe4qeoScfmYzG0kF4
iKmYMJsPnYP4lLtdZJ0llSh2aQqzo5ogJEDDpKTkhsU5n+CirU9AmKqfw8YdiTznL7RHy0dEae/R
h00S1Y3N92vkdEMl3tLiAHA0wbqoitDwagwG/OivvzAR2mFVovzGNRWOrgqgqWwLFvD1g+3w+71l
w2waiu0TKCZnIN0dgRrCHqjJ2Xgd5x+E9d1JNMYF8HU42JD1kUIaH6Ga4B3P04+qhfHL/ZP6ZqmL
r2cXaq23Wai1Xq/vUd7ZoHzMuSqUxGUusXe7CS8S3pQCTHR/4a81LUUHgUchBMLNAHnhQU9JjyXD
469VQJgPDP7ECNn3aO1HxReenKl2U+vHSHXDVK152bFIofGA+hrXvnNC4Ob9Ro3x4zo1/VxbTNCp
vO4nDqLszKGFiYnEIVVeg5+j2M/9tGZxdPEO5uA2vCwwn6vafDkZcRWT/Mi0cH8vw2HnsDc6IDv4
IV6G65xoJCSqA2WpY8w8ozqm89Rd3vCLEBB6MGwzDCUbZbb77GHRAPbRAIZ9Ige6V/QV1pRfv0AF
yOWmHg96GkhhZkyi/QDlxFVMg5466DlfcC9rU/ra/jienkpkNIk2lH1+J0InvTTR+IJ0lLShDTDD
u5wUNIz6KGVcqM9GXeFEi3/AlSPzWsluYVu6sQBDp8s2lfbnDy0QihhwoPQ/J4mZnJcWOaw9qTtr
cai/T/QKGhuXuSg+p7Dj5dyIKitym94BTrxzCgHGY1bONLgikcPbTJWPOzbAsE+um9Pbh1kqT+G/
hX0wKXTzxDxsIgfv8M/2ZHIAeWezYWO6Rf5efKEQiJeHFbQ3/67C6o3AhzQsRNQ4CKPh8yOTVEm9
K1Yal6/jZ1OPld6mo9wuxHgWRppdrs5veflJxLZlDW4V1aCM+3rETdErcK3BJH/Yk93/R32iUJeW
q6DE7BaUY82dEXRHm0VKDC96WiSOQLNDH4+kxv7eA9BN5WLIPFQJcOHZ5U+QgZXjn9R83JtAI4Wg
KqFEdYURHdYMXxjAFqa2PUbnwoR4lN3zW4hzjM51jxUOszBsUESBzZQ5jhN8n7InPvxpPfJuK8TM
/W1I5h25fzdIaIHYYTa/6R1pSZYnyuioiLgwsgjEaouz6pFvLkyHmFls910fhF3yQrxxGQiIElAB
TzcgdsS5WitTJNBqwRj83u2YYATK9RaWEpdRp9axNVqXIPu4I28n1+oFWt2DN8v/eWKLbMwPKbXN
ECoNKiAZYkFD7M90jAPRQ5vu+9hYKD/Dr6HA/OFkCluH+lzcwtji5yL3KT6r6EGnRRjD1JIEf75p
mx2h/D536oEow5ja6DosQieTcWFOfmd0DJNhnbUTNLV3UyFIo4SKk9IPGpfYb+z1ErPu626tzGft
6LJ7QgyNW9hehymGtGyw6CwNOh7HUb+pCKTK4YujW5hgRlNAm6kLJeu+BP6etWIbSVz74qnw204H
efwyXkKdJyiIbE5bdq2Mb0/azYzAPTwWkQvBMtgKnULQJFjEhfRjH8/8mFIdXftDY1C+QCwRPK+g
9aU7Fw7iCZ8BQXCAimsI/9/2efCuKFT7NDl6z45AQHoN16wtBSDtrcpmUqh88/xHLZvRzN8h8BjL
ZxOlpnliOJGkyI7KIFCmikv0IUkgCEYg2ouIbPVraOgH+VBsrS2GUpb/jrY5fLuJgCc9PBN8RaPa
yr05aMqveNe3oI9Ltn4pSQ+F/ujw/EfKZlOGt/wyn+Kzk6AHi5ld5CCEscwT+bI6Vm9v+Osh8PSD
iL6aIyZIPpNtFtSu102wcKNMF6ApPTrIB4qs4jxhA3c1Po3HD+PK1qIigOsyMNUfvDT2XwW5Fz/q
sO8ShwMSUoNB7zwYWsbbm0QlqPcMRohlRlkEcB+AFnDHbDsgDxDxsZQcXJrCDnoitIFsR1pkYB7D
JozVZrJYbWRUgPtwtRX36IGLaGddkePTjnf477V7/nD4or+cJ8jOLqldbO2TL9TnYYFgkw2eFeta
l5rreagwqGfYrgRu/xN9ng26XIzRGe6F7+bAJQ5DwpSA5E/2o/OAC/gM0RErGd0mmGGBt4dhDExx
WddMiNhGAeKnVN94B9BunfDwnorV+9O/Hnw5PkXD2xdaFobzTp7poN8eSNgwQGSbTJ8x3lqs5hC7
vJOYju9GkqDIISKKwzOZD9vmdx0sEVvPvt5yBsJSdi0sSI63V6js7jIfBBDRZUJS7+HxW9SX25n+
c+pmoAzx4fOKF0vEUcZlU+WY2GR9gZaSPS8dYdZjaSXm8PnFgW28mois84wbkPEnDwY6w/jnjYBg
Ev/9+MxrLbndt7Cvm7jW5IlmlduIlBr/QRrlQb2eI3udd4e3shmka4rAtY1KqFz9+fOdWvvaBS3V
Unm9rWdQs4DCUFIJzelnyWO7WrxX968PLHiM5arb+QdQYrz7dAIkat/s1YwjuytRKbUlsSF1qSkG
r/9VIxf6WRrpD0RJT3MxFQS9tk88u0spzVS9Of+V7Uh3W828kzoFmXfoPIp77AnzzagMk5Dm6ik3
HLVnkWdFGtHGt7s7iYIfD69tsoHe5XijXP1FBtfu87yrFaJWjyQDNkvl5UFMl+IrQYifskgixvmT
urXCDKGgf9lvlyNrUNLB5Vr4GCKrrMsExpIalM62r2Z2ETVctQcX0y2fqPsk9vDroqLQMM4nY2kI
0K4D7CpbIzRITpGGeaRooZdv0Dnwt/BvtkMjio7TT4WfDYlVFjP404WUHA2B9L5itDdeDwly/NlI
GR3nupDzlG1iJGVmqo15abdXPF4jHq8s7e8Zza7iIZkNUBHo7cKBAPIeJEoOYR7QU+iFI1FXcLvH
WoEGAQPEFw/5CO293+rgH9mZjdBNIHW02N/aUQW2dFX2yP3H5lnVWQtSSysC08dPcANNKpX/CL9D
wW2mGgDld+xnBgTFF/YLwM3OWYeo/pOA8DMZhOgQFFuaQ4jAS7/zM9rzRDgkCBkI5yOId17MMD0T
KdI50QBpyAQXKlD0ws+3yJFCOqUSAnSmoopmqRnx7a2aDqz0RXtDB3o0GedwYUyYiMBz5nYtVSE4
BfStC48MT5S0KzN1agEXs19Ul37YzMSU7q/+QVOfl0zRBSGxPnJV89H1VQtaPbFKX1j/rj9xhQ/1
zVFAZdlpXiOS175xX8+3OimU174aSNqFYICBXCPcLlKR5uSmtLHDHCXsxTsxWXJ1YkFHoFP/8jaB
wQeGF2PGGmyJQozZFsEa2uVO0t/0D0RZ3JLDfBgMw8Tf/DPR0+gPy6RmGvqzvlfEYd/ohLpk7e/3
NCqSBrF0PXIvQ0LIHUxbZe4ikFLQa4lnNvf7uBbbHInsTPKwJ5vhc2XpTEUx+2HrjK4cKvRLTv/f
ihl5zzfsMJf1vmw6AGXivYPjkqrIYLUlP1c8/Mz+AvpAaZ8BwFzNkELI/Xe5XAZwC5qTS4azgXzV
JTDpBYDqisTo0SgVClM4oskak27nOA02UjihWrl83VUumzq40zs7vltawGyJdD+1+CrLqsdO5/nB
Fh/aljVkOLHM3E2cwAM73UOeOLt4yS4YPdB9QGllq7kc1LxbHthAc+Qk69Eq13oh0q8fvohoyNTb
zx7XHEnLQx6GVNPSPetH511lHpyAeB7uL851X8WRpqL4H8JB0Lhdat5aRiHKa0KaoJAHqlW4aoER
TW60lW+2xcsN4oekG1p1OGEX5jj6gHkPtQK1d/hIQ8nmCJRwek5XKlAkCz6YHbYGqksvTlMiebg/
od2MGlkUYvZKm+P0iOC7OS8sT53Cvd4QhXMlElGLd1tfflOEyryqLkHO8VpsaG0FGbwqAkdmCjHc
+FUit/0WTj3SieHMaHVS7jaZPTkeu7DA+oQ0X/PMtKcGD34DkOgQWe0bXpjOp/33NsThX3jfWGcB
HDHFyCax8TlRE7USljCsZJow4m/HWkhszW2CnrohCAli2zz7BF5rY4c7YQmzmRnH2tiIJejrXvr9
mjnN1+jGSdHf2ZF25TbRSktyMVTi3tlTvyr05SrSFEzpqTijC/BUUegdRSSDIEbaKPQIx3YNDkRW
3FZK/wm3ux8m4nvHMECgWe5qf5OgdKkjPnFEwkcafR87YM67TZxapIVxmQSkgFfRxgljS4dI4KGF
FIicz0fQX9iTHVOmrcpc+iDZ6sSmlVGbw0z77zZHdDUmfuyhNpcr9GY20BwPx5rbmHWFwifFQYr4
wc1JuUtsunQSjqLUKDagwF+bkyiC/g01F85N+RZD9NxofLVn3R2Nia/yAVitwEIw5ZsEY6JiWKZ3
48JMY+3wjzFDYcV47Spd3Aiv/Zy7VFN0Ddl41J+/ldIVoaXleqA8Paw3nGbahP07dtWAFcD2uiqx
hD9sdwWnM08JjsMJvNE9XZ2t/lqdy9UDUlXiuO0h5gmGwpWjeZ7qe1IhCLZAlsnekdhJZX/46xBZ
kG4n6wq+6Wx/xATC5ej+T42oPknHrvmNAKeQP4pCNhBAUxQtehomf+Aiz25A9u6QvDXll4dCobq/
EWeYsdoMIACfMv7yc2JLeFaAm+AdsTMKy8N6R91shqTJtkt7RS1/RDBZPyAYb1GzWWENQ4V3PCda
lyjvLzaeZTa3dqS6sGSweEDJf7/NK3pgLc3bHsRlGJ8h9YUhK2j2lG6cgZ7GYSE7EwW7fv2IaXx9
NLJFlcjab2ofSHEQlAcUlw/WA95miO5vc2INXKVroW3WsDDqr/F4D+h9GCJgk+Jel37iQP9r10Db
oNkFLi4Rk9/djEUobf7gUqIWpu54silu+qlnMCo3157KeCxfhzkMtjzeRWzhJq9lYOO9QwVP8BOn
3Uq7sQ5KjHnpz+Qj6na5n11zDo0PaCAd9rkJhCyG0KqT+8AKpGBbMWFScfOQjenzqu4v717U17Hu
SADbNuj/iXen7FMIp03Jn7KG6W8xuZWtpIw4f9g69ZPG2hh9/WsTINsCBcB6PCxRiArjCG6u0kNE
3V4EhiVdSQRON24QxWb7zV0TB5IZ0I9NBmGqCmwcNR7/JHme9Zspiss3uGsMIMMcPZWCGoHas4uc
1rXenLzZr6diok/UZpTGsTfvgg3YS0+Qd5k1GY3hqRUhOYUYoa0rermA6aZ4FEQCvIO9ptArzqmL
lkRdWu5l1X737S7aXnhuJz/GxyEGxGUf4h2s2wpA6QDEmyT+LoRpnipz/4ttLz9yuV/jSK0gBee6
nzwxLO2/n3TbMcLHC4k1q1JB1SYua3EWZ1xGsDO30QANhfwDoFNTy+4trNz8jH1Q69zY1hS/JWNx
X4l57xB7K4iyhIgMW6s5nCJNRmHUcib86ISAknPmTk7RIYZYKV2o4S3ddAbn3rd3opPJV+L2PNpk
hXSXlOgzPEuZTlA7iVDg7CHfkRdMyNtjqEcF0iGD5KmyX2s52hwr0nXzsxFAQi1TtgVN2imDBm20
FpERCcyD3bU8IWxBZ3mScxxsk++TkQlj5SjOZpi/L4AlkTdkhWl6i8NAr21FUOoJ7GzEbI4qGbIT
97gClWKn/s2uWutLwoSE47r+ATQ2zHxBLQkwlv9mA8VyRC/jjM+h3tR6t/989WbhpDmfccbSD7Jm
TnoGKT1keo5ndG4ju1Pzxpj7bIHvGloZH+yV7xijF+oi3+gbUF52ji4XCQxucQ8vBMkiFsKFgPgx
yssrt0YeLZRnXh3MFTjnI+uX8v/Ars81S5cuTHkpBWFhr5So6NMWooncq0F4XvnK/fiXVI9vSvVk
6NgSN1U6DQV7opMqCpBHdc38LxZ/ZPOP9y3WPNcWCev24AWBA0g+LbW99K40vQgu2+CgUxKxu5GR
FQST4jYYUCz2KJl4PcV/zhfc3szSZS8nbB2INy4rpo/xmVhHx1cl6AA9NqtVhT5Bi2hBtzV+hUPX
+PHg+wo6FdfmI3tjKM3e8IfRhBfLggGCY2PJfK3KgEcqywvBdvQu0+pG1JZlaGNsi98Wf5rbV93Q
sH0HTbwFB6gZ4nuf3RY+D2IB4UoLFFaAunXny9QVo6+js1gu/S4cXnOKU0AsfAj0ORdWgVACkaRG
XrhptoZ3uVejEwPXzSYVyLw5xyQgAQ2tYTDrq0Rzgs35Ym0h4IteXfhU+qx2q9CscVK6rWY7nncU
jYCSzA0b6dMejYFS5iS5xRXzRB4I6N0rchkahV7Tj8M0RWZ8n7u82a8cNMndgWDJLWg5HRr0DovW
6ChhL1Wp/v8X539JIyic1HaTsHlTjH/gI5olzUrWb+5THGZriL5YG8H+JFohTwMwtz6Twj+Lrs2f
Mtb2QiyyXOaNwQpL0Nx5gil/Z8y7+cL0xcEI/YEtCmCQudrA7U5siBj8Z+eQTYBd2CIno8XY7TWj
VxO1Mrb9MGHn8APila+kdEWPqk4BiopnFYIk4ugUFU9M8rNlDzbaUKM07Y0M8SJfMS4nOr1XGzS3
9C6jSUsJGHoWHam8M81u+uUZQ0N1Vfb/kYyHy52thibUGXVj3NcnZoZWvyEtBoEDK7F1T7vQVhX2
nFFUyr6grj+xF8qXmgcBZ1uPVbZRmPY6WDFkYLUyKG1kZXfkhIVlwhM5l5h/hhwC62Vz/7pj6A9p
Zv+9KQ8jFsYi26dX/B6e7eO9F+zYhgLVAGakZwXUVf7XblfDbxgs+KkOX/0PG2rug7X8LpEqGMQs
rt60cwR3y28wa+2bIgXYACgIqbwmz+K26ym+YHgx/TVgIl/BVVS4cUShse8DyGB11WjwtPhnt6RS
35Hg8rpIQtf95yIrsEyRDToqcFBufxxtajUpuAryQYex+4mU3jqYUrkHHCxX1t0S5kX8f7B/h3Zj
BG44c2cC3SBrtyE8zwIa4XW1Fjdlw2HDqFaA3hNU80aNEPjWthmQy/9GGCdAYhep7//RGZ7iDz72
cEBy15kAss9Zv6ExonylY4gwc0PARRZWG4jmH8W6X6t9aluJBHQKuyoS4NoZ5useTOQasIy79vlu
qGUJ21Xm7Bcf2Y/RVneFiKyUwAwF/pvyqjgQQiVjUxWzFyoqi5KAVPJeBeUWbgSlZn74CsD1d01s
ARcqY92jZApHEXw+pBra7hxyAFZLsHETtIjmkF10c2GN+hcwf9EjQee+c/KS0JCOj5h92oN1GG51
AeLqwHlk6ZA5gOs46ErtCNygo4BXacRLQcv9wW3OyCsH3SgywTlcqFfJpRTUE4moKeMzmj6h+jEJ
qUts6f7V917X9pa9NjwUReMkYfDD4zE4U86PGs8x2vpyOiUCXtV/AnuKAPsZL1eKQycD+2jgi3Et
o3cmmh/K+5KItQKsd0CYB6eN3gpQtZ23+J7XnMrcblf3A1NVROoJsezo9nb6QRGt9IRHXU5q7XQk
Bw+VoBR7BZDwsvZl84Ccrrw6S6kjJ4bUIMGaTgUpBp4G37F7bCO6oi05pU5lB6O2nz9sYtH61eW+
GifKJblQBIT0nNEEk5A+6M0VjHeU74Ccanw1ss+94ymV1N2QsS3xUNd3Uq4XQltcnI/PNhMIhb5D
NfdpvoAaxew/D04trxZ9zeZ2FECC9srmAcoHZymW9MpZJYvzipXQsVl/3rOFTFFG9iTvkZmkDhTM
YiEXleZKgS2rKnf6ZueN8kaR7SkWR5WWm+7/sSU+B+thn/84WqIukquBANWMkjqXVoN3cP3+a8OR
B5pdQc9LQRjOlzfxyeMjscZ+WSteEB/YDEZETmhy5X58gBvWo1oXP4cXhJEwg9ey0jnxFLHn4CKw
Upz6bo2Q/pIsGXofF39w6Bai6E9HNODMFQYQXe7RA1kI2v/VeThATk8W8NJrQbXnMuThGJwAD29O
bALs9Bqai8k8zGkUKg212DiDnLlFzCE0YhdDzcgKDxZUfu99grDiVlvBGvwJxTpoMWg1Pn4EQxyB
QUkLA0nJRbhRukjUux+Rsou7LsKgOJgFjcuG+wK10xbxfxC9XapBndHiOe65HItn1i0kYURNQuN3
DZIjfKsvfxVzQKuFm0tO5e5KEfutB9Vn0VOadRRZyY/jIG8cgKF7sJVv2gx3dGC7UKM3L0kOSOnX
D/f4dm+ZSjEGp0uTHa2RKUkenKvB2FtILWJ7MLXtriqGakVS4wkSLmm0f1u6bCmTYlTUn3aASlL2
HDhWvE/n8nuSSujZNwc0M+6gZf+qSkL/WQq/yAs/Z4yThZAQr8XIYy5r24HjPwqRQjltzuCh+7eq
qoLxXNUSTEYK61isnb1wLQlTP15A80JB4lQH3Q4bQEQ4xl8umeJYDoe3Ie2Lq2CBmf8B6CrodVqO
Ybs0C30L4LoEU9m+ubyyagoW6g+CNUMCmEfUuHYOcjd2IzROgMzRJbXz2kVJZXbNB+webUQtgK27
PQI41Ly76mF45kGVW3dguw7jWrEqL00OO61x095WPbkhnhfH642IIK2wfhTNPTBtKLUxc3xgN2LP
qZOKK9ATtBo4PRDtpLmfwofDbJHYq7vqr8gvnwF53fK9XBfYzerv9JvCqxQTzBAW5nQc2mZbeV2v
bFnD9zzRcKHF0FEomSxIrAH3ghh6AqdZ80Lmb2bxPNcwqX2wckoSmD4cmoz3G3uvTTO5HMTPtVPU
H8Vf0YtNDEHmOmWXFbfRo6cNPCkX+Rz7a0T7W3PqCVHgBrSxnm883WX81+Y17YYbAxKKBgaBos/9
5nwdLCeeuEcidojkEUA8Hf3rx6s/RjfwrZb32aPkUX7RIcj8SdwmhEYLy+HIsSYBXdV7GfSUiIKJ
hOkJZuxjnOC/a539snVum8ylyMwDA+YtVs7E52oK7WeG/KoM8/Ixwsc7VT8r8Dko/OFyreOEPeVX
H7qbwMnZzT6mrbBBmkp1eMUCvNhkynHrr4/iWFRNJd/E2nIV9j62ak9NOWvjzudArCatumxzefZe
uY0nW9qnQliQSCjw50xRTwSHb/9mA2BGrDDHLn/uBhTKap3lmKlPaIZbjpZ0ec+puvzvLX7O+UkL
3FHRRsVucw5mQAA+IU4C/srRQLWwAFfKCv1Dnh4vFn2QNAOMmKgfTD1KFF5Kigxy3BNRwVYqrwHB
Q9XwTo+9tnfLuPZYZWc923yfDP9+gHNspiwRYzugscviwdeIZL8ruusl+rFyhFMiF/6xf8QA5DZA
JwGd+kQ8vVZcre6jXX8tXE1DgcNxZKM+HhmdL9AX6DSg72COoXYe+QVaFE5zlaG0c+2AviFOxiue
a82MC+sHJuEiBnPRIz7099oa1Wswug/6ovm7gboLyJVN8xPMP/aMB0SBmoBdwZK0OqK7rljJ83iU
lGwGKDQXrbM2ZFwuS9bspNdRcG7exUJt8VZRpmPF30yCg8L+3hOJhsIDJ/6V81KOvaRolBsC47Iw
TAv4Q8N6piPe6Qu6XD7BIXNVUONm+COiCXAYFRVt2in+wtcWJEFoKPG/j7gTjnypFQyhgjIIGoIE
xc/iXkpbheXwklQcbv4pRASNopBXOdbsZstETVdxgIMIYy7OuG+m+c/A3yqPQmxeg1UzjE1k32XC
0eHhkVa5F+Vg/1/cNMT4Z7HOBb7Hf1qsVfycVKuj+TK5bRGOiEcPUXRvOEcDJ6xdLYnW/qjj5dox
dcsUTuaZ0cg+IqPhd6gYe2GFqqB9btT7bVgEKmJhGvpKPJPwV0SiQ8dwpSUmwxUcztGPJjmMks6+
zLkp+XNJdDE5lormdnrN/HGk/86leU9ecRjKX7/b+ZseywdqLCTxr3/qJjQwtYWWIjt5fxci+jHY
ZILybepXuG2aAZA3c01RYJeq5DpRBlK3O7oKEWb3OOOMqlkLxpnFa2vMBqKY6BUXpwUzVSNmCxGP
cNRQsEJSN4PI7gfXvI5vprc0kjnBAd+Nsdj8hC0gf7jKA0FBm2xhOIT3aPaxGwJ69UihCouKotoQ
0HMZW0qptZPFmaXatn/NohpwBjJQyXFA9QAUAXAJTEJwEs+ga4ofGUN73r8ZUSsLrYqmyq3H3Gde
XUieLN90pA4CTk03c74ueIGa2QhtsHuRWO2ql+6oWll4XSXZ2BoAzl8TuxiNZwSLp5+/gA5LiNRi
O10PRT5LMwMRj7wLBjNcvBI+9xfkgjoOESeEqCbZuYziuNfa4lkRl85jD3ZuJGK/i9V+mpvHISHp
2x1QxWgRpNGgAvMD7OhL8oJcBTBH7AjtLjO2QOJH7S/qqONJZs38L5qTKOVDLt3ENi8INxK3hNUZ
UcH5rxwbVYPN7kyAJDHvX6TGnmODxzdww59IwB5khYIyagD37/5x2P73RWcAC1D5d/fw7Mk3+efX
hYaF9WkS6J1oQnPgQwgzdbrMQpJoB7Q5hMVdbYesPC+jqPtROAjA5Et3al7SMZNi3nrTobCo7fK+
jpap9q2+79mVC3BUsXWTN+iQ33x6QO6asYkSPnIAcQdYxPzXUMSSIXVJSm7CLKvAHNdqQjjRZVIz
eCUe0adCrX+z3bUfUtodXNvcaX9PZdGjUwkeltusN0V65iAuXSOJxOlqaEOQ+PS8U5HXqiMD4i4d
Eh8ul2Io4pQyRnUYlvtxVMXk7nKEPHsX1H5NcsyGDFAbJyou04QVYp4t6grUMhpzt/7WNRmPvhVc
Fleuv9ckzugyDgQtT/4jhGzgyxYoPuZ3bdSAZbzP8hwSJHCi9lbywmqDlJg7tsrVPqmPL6HZOkQl
i8XktAmmBrcK7eVa5QcdCizKGEfbfq5aRpJT77j3B0gh17Glbi1X6kUXQD1NX3dCApurvzU059H3
/WlEUn6FZprEDcngsEloBnHtke/AGIWh4fZ0jI7u4zXtBJl3yGWoUVpi6Tdg5xJUUt6ah4fZvW/9
7g6JRzFb5t/XRHgxHDrEg4BK5PBi80LVDfI9Ldd+uEX4PJp+E2cTv0S3Z393EKUEYs7hbQm57qek
EFUUXuJlX4lPOlnI887yWD0cf8LW3Dzu+OfTaqoTCjmkPPDEqFWv0bN13i52DKDg+nMg1nYsBPka
t0Fms4HZ5y1H8V0takXu2X/qyVFm5tnWCaPSrqLe3EymJu/0kkFbtS5/HN7I0MA1Yu0GfhNTCJCd
A2XXY0uNmUsZBxvdSb2XUEZtXhv8KftD6NvIrxmeZLFyyrzkO/4gYF4wiH12lP+xFNJ5xoNdXXY2
4NQv8Xj11Gt8b9ifk9B2Os+3lAwqyejIFCUCC7CycEzZClK1ccwNyogPOi6OskPj2Utw1r0gTbQ2
HgxV1Le0fxsjoadrWgCQcmr9M/WEGk3xl9upPm/jhddSlO34DVKgo4TWGKeUdj2c2i3pVxU9civY
9Y3XhrIAUCIUwFgkhxLDUE+spgKBgcN0/m3WNO8ZCJ627l0ioJUtGqc+jDgTDAVssFchwxW9Tpyb
gef1p3WmWKbYLhhVpF8I/H4+v+qDqCmJpc4pEWh7xBrbAY2ZtX2b46T+GVFXHNllXLkvbsgdSprh
a/Qg3gMmWHrphA0mBczI2e9gRIRa0DxksymIVQ2n+VhIBUMZObk4agdd1KvLfq0duppHqxBo4Fl5
f2CglOeGUc2fKYwbtw6J94fztqTImjTPruxLcPgvY7ZyrcvWOHn1pl/S/ATGfb4C7E9dvYW1Fr5E
yXzLQZ9uiZJ1Vn7E3j5NjpP+mknwcqjwmsCJVHuijzakVFrzZd9Sk05seg8IjJbN6FO2oOjXe3YQ
IvmKS8YN8T8SrVYidZLhnOgsIJIOCSsr39VKTk3w7Eh3JLszr0gxImTXny3JBGJvyP4Gy92N8YZd
XvWG7Pd+ADyDJJGTnMa7ysAJRlSlp0B+OXSuit4aYKIVdhZQmT9aAmKtRbb/vK9phgylf+pWqMXb
C2pjKTvbeAFEHt0SmAR381lU96pOFkxftAZ9oAK6AkAqJ3zQZE9ylb0cUn3QFxEP+vkEMYesmpv1
oz76BPOlBDksIptDs/OnJcyMcaKg2qbVriT4TtxpnkTpxnYT+j3NWssG+TGtXTvapQZldfNQkAZc
Ju6xZbThj9UFyWlBk6r3fjiHJ8kWCvAs39ewE7QfHDlagpOKDv1N+sSlOgQUNBHxEzB69+Ks5/3r
3Z8LMwuRmlJ2fccbngS/H3Gr25ywypUMt+ARJ3bqicmaKsntcP33zEgeJJXwiEjKKGZzhXEiHxOC
Uu6xevgmJJpgDTdlxgYycCF/C+8ervZBt3UFrpB4ztqf17RZXtMEP9y0TiBYxhDu2CAN39J2hhVY
312J3QEcf3fYT/aC7YgfFEGjWN4L0ixyGS17fKoFID6WVd+1PjlH4BdGaGis0Vf7n2BdtxK+1EIS
w7Gz75rTwVGVS6AvqUctMp/8BjdgQQCojmgVEEiwhU6CKNHruyhGOOs6MJsFuH4fH4IWR6s1P8Wa
4B5HcFUCm4yz7PMgvqT+lhCi000sp7+XnoF9LvS3NXMO9M2M//kaFCOXT2+JacsWkkj7qSndWXq0
fdoFXEmT/5KyZZA2+VeToGC8LZbzyX6E0OZHEP8mC2MFFiscx5LDO0nDkhFcnDLKHQ6YvIPfSu+x
DNW8at1E0URIvhuMsHD02Ru4Uyid/OUAWOYPq+JVPzXeug98X2VdsCS4p2a8yB/skPPKu/7OG58V
guKoMjhAckKHnGO/8mECsYR08iB3mX1JcXxpOxB5dYT8BbtmJJRvSJlnC+6HmMFo3GkbGlvlc/Rl
hYxQJe6y2ESl02/5D6Yt3MJLM5Lk028uLIHbDIjVbKyoxwjvht6Eh0PlKrwbDC75EK0huyzwUMrd
8CdPRX9x4iYsxgQHVLjLjnGQX72ESCawtz5B5GtZWxQxoUeB5INYRtQpGhDLDc2sHs+JpYDBNor3
G6adbvuc3ryCeT6c59pkf1A5jcK7BKN96l54dBu4lQvcK1nrUb3laAtuk5kOMOdIn/mYoHrhltWU
hb3LyPkOCRq3dKib3kM2RP/et429aYHnpIh2jjO3uQCOuTIhJyWjjKllTR9z+dWJbusssj0MebOG
2Qyg5+mDQ5xW3xq9j5tnArqHaLiXu9uMv61d/sDmANeZqd5083jMfb9B1fDrELdJvO/IIgMOA5CF
jAqxyy9fm8Qky/gKW2dJltDxckb5JBXU+HLHrE4gJfkZixfib5uAL+mt4NiniN4Qd0Shd4RaAC9b
6BI826DmrVgxoYQm3Juy0EWgS7j64DPLJ/w+c/ErPv3Si0kRKA+qCpVUalCKWedFKNey85xmXANV
ltz3ukvQOrk+K9WAucrmXS6gC7NUrkk9zg5r1IUzOBxyuZ1H3PCqE4Hbi9r+mkxmJjE97F9nNaKc
uZvtZBSDiMmviM5eQdKxqzyWsDzs5XcjaF0ZFE8arcU0RmvHwa0i9lXvqmtHgvjesUvPoKKoaLpy
bP0JzhS7NHqKovOu2FEjoddaszpL3geYh3ovD3EdCw2eHaNXqwg195oNTWrT5AwJM2PTryYnSJQJ
rV3x1qcfWbJBhMw1Iwu0OKkBwDQFOuN/XAeI5ioZ+jvwFhXpKZexrwOfA/Jmncx1KqkdxUw5xos2
vokDyiClSW8boNoG48wXIkbJXl8D+exAwY7nz6PV1WI+OeeaeXKs5CfpJTQvDwzqsYWJk0j7f243
gfJPezpUJRIsidgrNImlpzRmK/dEHMbzveiix/E5zpADbeJVZp5g3mC37VL5uqOy0TppLlGBTbgz
PuwA++pZ5CHRJcf5pmx4PyBAvmBFx7zXoDbpWic8qPykX2kZ6LgkFnP/RLmc3dd0A67loxiJ8bHY
27YW2ZVacc66y3ZK1a0fv3OgaWnAy2CTPiim/0Lh9jNPP+gc19fK1BlQ2q1PlBthBb/YDzLm4ViW
8Bkhh65ujdV28jqhAr18mSu2gvtSw2tV7muac0zjGFDNcmYyoFIio6kwb+NT6ggd9t8V8ODrFpR9
GJvOQYw4Z/nWJppVQFxK7XgWigKTNfAV0DCp/Ijo6R0oUEuyeZcAxH8/QAzpcLeZ5qoTzKGD/np2
m6KIhzivKCqo0h45zUVMHbbiNupQdqyOw1uaMfUDvOD44l4ycCTNVx7em2IAnaqLmp7VCu/60x6q
ujWAVq7tY5kfS9VeDNpfu9b3i4xluKxjbSszdGW+Ae2u9DWgQrBv1J8T62TOB0IyQkdksk1uShsY
AMtTdYxmPAqEw61r0uvafy2nCBpc20SOANzlw8cyRW1ny+CoGV22GYhq/Sfu9gFEUV12O+q3Em8k
ws8o8D4dLuurCqXWBx5O6Ne4ZCqfFl8r5HStBvHAyya9JDfXMJi9+rv/x5eEc71JFJuec9AJthF6
vP4tGn1PIZXXsH51VR9pIK4I1ULhEs2mrBGu+b/w20oDPCoYhq8vtcgl46Jw9d0KzQe0TuO70kAK
UO6IZSTZ7CAE0U7tOF60Tf/WwvMOtkXWUTobbIaF8/6WABwlODtaDYpKZqpofgyufJ6vWub9TOEo
85YCizv8OdfLuLqjZ/HsXVZaiJ6+iWYx9XmSqL07m8Y/tqZEoS7pTWQOc9Bt7EXPvAx81Q9nUBtl
+ZZj8MTwq5N966Aobtlhd+9XEUF4rlPWxHtKr4v0VxZm0yWW656oyZbf2NepqbWi04pmF/SWGOFj
IJt71tMMP0V+EBOmstJyYAxswPNjQ7R8yZONw8XEPNizZ9Wsc1dLwrSBGksU5rJ6qZ0LOwB2/zpY
RTuT42dGdso3oS/bvLQcjGyBp9lpKBMriPjfc93rAbJiB5F6wnMzh898N5t2K6Ajp/pQAalrOOpA
LQ0o2VIhAwu2HOirVkuM9ewbJ8O+B1o55NYR7TXtQdnrL1XkP1STEZQ18YEjbKhZmHvKrNrZDu9M
CFe/09bl26N0LYK8WnhWbxH5xyxetLoAD02JsyO+bHJDGmOk8UeJY85QfWMRqztn8vUGbqL9L4UV
de8nuLI/8LIuiVN6hPn1+j+4dIr5KMjMcKzJAemGHsql1NehAKefdJxNuUY+4df5BC3z/07g8A3w
p8hUqwwDB5YSIaK+S7PZv0LQUX7Klxzgh21VPGpMP0PYKFTX5UuumDgCOQx56HWU2RiQ8gKLA5Vn
f9SnYR3h5s337SRf1wzYET0O4aU5YZpgIyQLpRECJkeTqtvfai0NdrHV01CbxYjkZ1zsyqAJ0Olf
5DGNnjqiYDKg3qNeW5UaEynGuHeGZx7q7zFb5r3i8DdFRANyDA1WQZyHim29EvifbEdR8QbSrSH1
SJ6n3Tu1VU52fZSODlIZQtxss4d8cKm/1JSXZ00BE/zbA71wl8e0xYr3tV4hz5GQtMsg41EdKP06
l1IW9Y2L9ghrEG14/Xae4UsDFLA1nZ6pfNSSZSStU0y3L58a+AdrlNHFUItbg4N63yerbhZeMcny
0cDu2GGZj5MDRe6scmDcWWoaXvyxOeAA2+WGNRwde+fJpxIiMIXzti5Hqw3CbbVXVtHkFoGLYrhQ
rdvhbidtWf/ad/v8ffo02hMbX6blSoM/Yr4VH1QkGaPwfJjJWqk+IDhELykpjsNIf1Np5AYSC3+j
Z03z0CqRYf+6kvo6LaraPo13yt55RPt0BlNC7ke4AB00Awbkdm5lzStnk7PGhuK/6yHz9xlK9g8T
i64yYlSeo3KYEWJhvLmm7i1tqiW8Qe3Da53LaaDPhPKUISWepv3fL/xAOcwk4Bk4c55z5FaH6HcT
04uWFFR/9OOg/e3Ci7UyqIRQ1Zn7NyxItXHaEAlxfGhijUzcZPklwLbmsnGqs7JcE7zDroFiwQrF
mEFOTBMlyBiJTZMPXezg/hdJ8rGIGLBBPBqJUIorsFYqTQvs45szHLpq4DrUUT5Hy28IVX+pirr2
wYtzwguoDS9dbjZuzUCVXs4pGg70XDcdD/KJfg6VJp2U58mk2Li/NDJbzqk90cmsQNQfNBW64eRS
JvQvqfIlNYmm3tRJhYQ+d+VjXy3ZdigXIbBOn5DuHLS0ThfcvuJe6V/tMK6o4MJrwI0CNyTTef7+
TTkj7JTt0WrVbc/NLQetBopo9IxAJ5kdK2nK+T4L2Bte3MEILXcgDBU7D+xWh9wrt9N/07j8m8Zp
YlGGwGOD4XLgiGKdmDgFoO0nv8fqP/lzG40R3o+ppaVvFEU8qVGqfzrr/KMXL1oMqaSs3eGK425X
R51elkzvi+95Eg+rA61mVHJtdv8qpypAKXMuqEgNHen0ebFewSod90ZfQw5JmqpqizP4RRLRHsYu
Vvrgq1Uv3m/KAg60oJYU0iB73xjfO2n28A0WoHr9qmDRZAgdo65wCiq0CBAWZpq9sw0nDF6xcvjJ
rAP9w7EQ1Q8IiTcUDKPUDQGTBISA9uc6eMU6iOly2YBKv0MDf82qVIDCvtn3fuVGkuyHIySGWBGP
2BM/V+0rcslBFvR1pokUEdlHGZ1H+ttTwOb9Ada/BZxeIcpe1y+QOMxhPu4MpfG79j1MLCBc/OFB
HuBNsEbuKW7HrRrK2seI5UL0i6iyNFU5YHDB6jl6POhPvudEXhqzpptgnCKFS7mWo8Vi3NNS7hXY
cxHuJjcGK3g4z3lDPEpBzmD75CEHZ1Yc1LSYtPql+b14xSZDT5Gh5aJJOhTJ7/gvURsrXLHO3obE
yamGU6O2ovJOFIkkUCZkWYioSKrOs6nTsxzsWt4XjadtKhLxEzDn9Mf4iiMBmDV8QYttJwX+Uihv
8tKc3fA7YxulYqddmOjjiDG0Px0Vqa7Wfn4YfoL/PuqYe7qEhndhPDf7rLRroftiqWamN2fKab/4
SbVAdW9l6P2mPpdvYC+yY3fEGdpHy7msO5HFZR60SqvOmBVo403p+q3PSWA+hM8pJwchqKbAI0n0
DzPCfGqXrAeX49ptiNdbPeUth24Th0G3g15wWsoy/GH4Zv/RT6i7i9eNZZMO+sLLqt+KlmzypD3d
CpTWJQz9SLzkvbXhbQgh/33bi/iGcupPcgYvhYzB+KCYWT6ON6ElVd0KqojMkZNG7BvYJ8zagYwO
kykrNvKMVXBPOBIABp3HrfiV1np1MoG0lmgfAYe/NpdJyC8l8MCHw+NM59YYbt8qDXaNfrqIkMcN
qqG1uFVyRd/Ruy7l1LLv4NKexDFLdOljIMpGOdJNOIaSGfi+akcWcg3q3OIcP9JzOo+eV3q95i1i
5pUUhPjSyVOREfCfzpFkHRbGl3FfiYO+Kdw38lZB9kWL6v25HR0Qvc8NQGOw62KvOiU8sShvzpRn
awfSzJ1D7SXy5eFNXVcLMoV5laqAEbzPBIkM7aHM2CNux7I1Jwgo1ObQ1yT3ZprVts5tJfZyiWee
wHGFuxMbG1x1VSqI4fyyWC7jaTzdk0V9GCZAWgXSZgg+ZU4Lc6lz3HA4p35KIjEDkOhRZ+bGh5YC
b6FUvDgbWcidnVG6I4FcVchP9nmksBz53aAd03qmD4wZlgyitZHrZ43MYq7A+8gyMVSEFYjuGNSk
R2ZRhYceD00RE/deADC+s9hQfV6bvi+wM8M220m5VPTcmINS6XDgN+22LBYu4toKRTR6LVyVG/aT
BUrD/oYmEr/E1LKHoz2RZJpxUqA2UGAvfd6yaTC9Mnq9OckFoq2lGVk+KBd6OvOPJZllWUMXkCgJ
hDDHwpz0PYS2B6fjm7eNsYjiyOULy9XraQd0/MO0AmLjiqPdeW9BAVe6++ED6YVKhVfheYNLy1F8
E+9v7GVQzIAo+GCztC/6m8ve6rZqEcricvaGUNesuNN6u5sjkvMgn8MhkNdcvyu6APFogpJ96GhG
ffdeImXpdNS08GetG2BcQIt20ZrO2cmQeBORV1cbwDmKa3cnxrIqSHHy6EeBcmkuH7O6pll+OSMS
kz/5xPG1TG13vlqzJLREaLHdFrKWmoVEGwmW52b3FabFzttGUmRiW2sytNQK+UFP6IOI+rNEms8J
lH0bw9BW4dFhtlPpFv3JrqPHaIUw5WXhyjZDCd+LrOTN6avV/imkmrzZzazaUZz4kuo4cdQgKY1k
RuODGP6tV5fysenpSNsbs/cQXQXiQjUmElN0jmuWQF/8HHeq6DVJXEOPfwBgRS704Rdjpr0aMOwl
AFOit5m2LZ0cg7JdhGEJ2p2sMQl1775/OaLiPG3HymMXxiJpO291swQqHhB7ML+p8YRQZGV1h8sh
nCL3i3gcP9WiCPwI+huHCCB1J7z4wujqOB98CM71rHD6M0jxzoOI/y5c8Y6VckP6zbscGx7/uA0l
YPqfdpupij+c8ApUO8YLsxgA5wDYk0lEHSLWKiiAUR3Tc0cbkzXmBmMqQX1tc1x8ADN/qDn7xAo/
zCncKj/Nn371dyT8Sx5VAmho4HEDDia4TRaOui0381bkDhiJtF3CZHGFFY1wVJYK2NeyxdMNIu2O
mOTwt/PFSbDIl7bG3vT/egC+JqxGks6t5CUM9ZoFP3n3C4BIsRn8v4hrAJaCn216JC8WWBGbWUqO
yPoSLZIG21nW2aZ4xpvqyiba9fvYUWkOhDOOWyotD/7Tlbb3r34KoK9TwxRvE3mPX4KwWxMb2OGI
aLN72MImdZgPZBbuydfyYuS8ftXwSFLRUqacJEDa2OrEzWDjqDII2q61kBNxRXFgy93yNgaHbzGC
Q/CigUnYnqkC5IB84wb5YGbeoDM58ZISzm0AXIdATG/tzxQu+7DQ65zxcuY9d4C4wiHt/bF111nL
AHHkO55riZ7L1eOskveVxdQGMZeUiBr9Id+nS1AJ1dcPZePlCGvEwrRY+0LNdE+CHBqON64FU8Af
ZcoQhHdgKCpjKrrKeM/caCUCKVivwE+M2wHJMIm5gPfiChiByvzmXcfug81NblAg4xW/Elept8CM
IGjRuhUo2u/S07qKJ5mm/nvTX05wvchLk5Nt633IPEmJ/db8WY0g2eZkOBBkXOVll51+fDdV+4jd
sn7wyaKKwd1Tq5e/lPeIf7d2wv/07sYFKuWVO5xCaNoT32JBMKS0ehRYgnvnHwnPbXZXvB/jZcPx
iiW6C8xkTK7AxMy/D8wN6ZO01hYolKJdFdQgfdYFULp0primYXYQRMo0IxMZC/3St2Z6TxvE+QPR
ovoYbHQ1ft3o0Y12wrMIUkcLXPxxtxOgdpwSk+84vLv3Wun0IXhWk6s1cCqD8lC5y9iTtjRlePE4
APiO64R5fLEVjbIKlapee6oyIV2fjtqHFriNJrsLKmblbE1D/jInFHbAiYEa5By717Rbu3Bgli5K
NU14Mxad/qBcRkftxuY84f2IER/4fLqqgKA5420RiwkK00V7yudehrzPBV6CAMBM1w2x6GwdYupw
O/6tC2v/a4AuSbPpH+yxRCrCMJfoGOXMx8xkZeQTv36Qe4eeCw+oA/yNGDQVOXt0aCzxTHmSUmZC
F3Zn7TX0BFFQBQhp600ZwENRabkJ+kk/v0FPnL0W8z1CnzflXmxxmg10M5W7nN9b/vXlggBrWc+g
mzMaHvNN3TOlaMHf3hgUIC1csyztjx7XML/JMS5hwjHQ9a8waWD3ylFVecQ1QTrFZKI9obsULin8
4uMI+U5oa8b+P/HG2IdjfrLzooHHSotl7LYHOJ2kB78DZx/uLfx9o9kJEy4Tzzz89AxW7g3qeojr
fdIkHL3JLOrQc7gP65+sysBLTDKOCHT6iwK14KQplisvSXJ1mhMPnEscYl3Om7NsSWa1QAd9GJZi
+ujBbIkk9txxJWp7EtG1eUJWpPR9ZM3hHiFtQAkukZ/yV0elVdJIlEBONy8vIK7vjfniph879E6E
HJlqXCcnTW4m/TqRcm7oJMaKF5UCJPARrkplxs7sraX8zRZaOWLyCV2OF93+ExnRfl9cuyo/GH2L
cyuJ8waRPk2EuXx3s28xsxxqDTkJq9VSmYc22bMtuvVRdQ/GcoS4lAJ2bGMKYACONaA7/FSgfZ74
IszFScf/AHNFhzutMsL4AfvR4i0L59xltRQJELeMeN4W46mv4VkiHG5njk6XovBOMWqykhQKCgCd
NWXYMhmAg186Zl21v28X5K8OtKNiXSuWEG8/L4E1kke86ltLtcWdG04tnDaC14sT5S52jDEgcZ1I
0dJImpIjsjN4Sf2dCZraW4SqMtcSP/+Vm1hFjbouLEwNyNGYhIELFn3vvkMFW8l8t4YTj4wW09LH
+UUCBm3y4/jwzrXOWzXtnZW6dGQ4wU2qYX+KWaU3AKO6QvW9GMbDhOdKpjfMRQpWPbn8HBMcpcOa
yuDWv1P0M8SOoAgCJ7b5l/F/9k+lqlQOwdVbswiOIDhp1ovws2hc8K7LSVPXz4k71qo3EnEXdezN
1kqLDcD2wgjiQ3WCvGYYQg/oAf/NnjkSGJ87GcYa3zBe7M88F8m8jQjZYamqryH0KeCYSIkutim8
5I6B8AtKUSTHK4GsRh3nb0Y3xUIrWj6TPq7GnyuzM+5kTyvnm4WVR372L12hP1z4Q/G/1/88PVIR
DsSdO2ugoQ7eTxL8DKSC1Gw0wMalb0Iyzjk5t11p+pPftpzIrJsY/rbLPlKdxUAQcpeJt9E59x/I
YCjjifBAr1JB1xap277dgq+g5CjWd59397PTr4wvL6YOEDWVBKdd7CogdTjrgt3jeH8419O0cAo9
WBXDdajRVWc7dn0Q3kHw1fshitW0okRAlHBe4Vf3Qa++OV0EzHh2HEYyAb37J4OyXmeL/kuln4/d
IfiM/YjQLjRkPKLFVRp817IwLj0/l4vnHQCe3tmHE7X/Lgi4OMeSMFiAlA+7ohdLOoVMJ6Gary2L
riKQhc5fSR9rVPnhoNBZ+6hcu75wB6KT6MHCWJKnuarOTTo8u668bI3/D2NwrXYuPRIOanyM2hFg
XAyJCIqN/vbP9E9owwZPFNnbRZl5Sa+KaCIT3ZuYf2+Fw8lHajYiabEbP6IqXM3xosrMlo78buh/
f2C6YeDVrh6Hj9yaJzhwozFMXoRrLwt6nHkgISgLYMfQ0tEj+xpKYgkRJ5DJr46wHOr1X51sGW1O
5HCxomFIthmkDG7mGOn6q87y6Cgz9m0/uLqxkfLn67q8LcYlPSHSTX+TEJL+nwyS1tTxRdKZdML+
ZTqc9F9neQIPVCmHwUXejfSjdfAPCLwXvwXYIASqZfQJp2+BSka6I75c4UT4N6+C+YyU7sikSCvw
ZuYkr05xnWgQ2SA7+sygd6TQrb1XL/4B5QoVneYDxH2PEcv081UHHzc7e2ds6woMI/0Pa3CMRFrz
vs145rEVahCF8oK7dPU+8NMRPJR+W3XDBO5Jw9l5LgQaywh/GC0HX+goAEP36GMelXW+Gng+udbB
IIseupVnO7rvZVTD6KmQI4vVFsjcK63m743dCv9K0yvR8k8KX4jhax9w5SCZZ/E2+Qn0qJ2FiVRQ
CwnpX3nBObBT0qLlkJuMybC0K8r/s2dga2ukgx/9fQ1MIg9DmZv2YtOnR84m9HyhfSqh+KgTpw4a
V0k/Mt/BMOZxJbZ+6aZaBESmeVJnCf2NJjCojmuOv6LlolsFrGpLDHD5ugFlK1VB9+78la75J1g8
WbW4KozPDrr/MQuaUvEvzSTINQIJcPeiukr2Magb8Xma3mzwFMNibshsBu2iD+/HLdz1dFpY4jaz
4EJ0P2+LRL9MBn58a/ahyw8uVZuyZgveSy6ACj+x9DtOr4DhY2o3vmejA86kvcewdmXpWmA7O2hQ
4su1vmjcGW0UzHI1H6TWpuiGiU3TM0ZncLJPlzXL82hCWvRpoAfNNoSJqt4c09w9OgoEjPJrbJ2O
n2tH5jE/0NxQ2RANLDTxfrKIXZMCygduRs7PPparFBmT6FK+xzQmwRsHZW8fRdygSsMtgAEzlL2M
NKe6kE2Cc0JtQ2ghUnWLZZWRBgVyPaw3qonhZp31MpSFe3hMCwc7IqNaLE7jQx6LM8PAVUhDnc5P
czLPOIDGXa8LtzOCcpZ0aW/G+XZ86XLMZHoyzBlnyxwx6JRudps6YbyOgt6PCW/vszARKi5BBBtB
4Dc9yWQgxAqWuXcG7q85VhFm85SlsPs2A8ZXyDraisVUK2Wok2oyv7u3B3Xl9vtXBDCnwovuXc+X
eYYBL0586gKkH2OeLrPPuk88zFonwZQ9UFun1OUPtVVnQ9ecUms9u1IkdFcZ5YmpVvaHBaB4s0+O
uuIFjvyyMgC5bS4KFoPXC6V7fg4pFpIzPO7dnl9bngfqhJXfslUzaL8FNBUGIYZupMRCokDim84r
NIRRWViEs7LxAS6o1J2yYjmBrkVz4erMhu9egkzIJ9T1mxbBThVsGmwpM1pC9yw/RPDhRUw74oCe
E/ze5zUQmJiPOGnFxRvyzsf8MUhZLeSBxXKGe9C9zlwzIaFcGhjeCTSoR6L9M4wwPaJiBbNtcbhF
6as8l42LnFlG3ukHnW6X9C2Tf3lPXsV56ZLdJdQiFA/b+qVmpwk/T8qC/+GZBx5oz1quTDBxnsEY
MwRYnaAEG8RAyZqjs3XM79NhK3pdndtYFfhnj8gXH3BcJkA5m9earxlpZnJ4APUOJmPMuI7nUIgI
vt+SavH1FD9hOYf1vQ31oYsTab9h8YmBAWt9Y8+Pp9QKGtJLh+QKvq9gHJpvwF1Ksr/xA15pkwMu
eCIQODap6XiXVobXE7/zltFNqwyetM8gqbz7m54kZ6SQjlLVkiE+/XrH+qIsnhIL3RHJfxIxaGFA
x/C0EsyDbVSYXDOsZAhST0qUy30eCC/PS+oHW+Zr8lJiGgpA5jTx0jnTxhr6E6Q3ChDRrJDOogVe
BcIdhc7Y0tiFoIwIPqRa2Cx8Qo4JFYgiUn7AUIbGkWfy/WwMSZsAHyqTsmwgCj6cm/1XKfhs+dX0
EDcLRju6fCwhz6LcPBcXzDqecxaAP4dPcLd7gS9ubGHTp7QExs84WV4v/wup7lpYf0+z9J9sCDuy
xc1y5MOMznKrJW8JX/0+zrkmtgL3tJVSLtsz1jNIQdKnZqSaFQ/pERGkBy+8/jtw8pRvEWZq3l2r
EgXIRQW65HAq/7bskueOS+53ed1O6glCPbC/UaD0tZoL3HYr+qWcvXla6lSHRv46PJtMz2DsloGi
PMHI80wnlO/3Gwm21fcsFBX1zAAxMfWkzHDL5hLfPuW4h/0EhBHyKxZpAJmD+yD5TVnDEf7MCQNT
5RX9bTxtXF7V8ug4fcLvR1eoIKKn/3/BfnMXojM7NWjtuUTzcGKchFF4WW5dxhlH013JGOiz/y2G
mhsJYYxbY4xudwHN+bkv3VxnVFym/L5lfcNfs9u+xtcH5epZ0WfkQ52XXwwZtRd0UMTw8cRtUJ+X
HPEXwQlOW5GMtPFYr3deTcBKBpzMSbBMZoTuXfN73v54vCOxsTCNGmETJUrWosN6bBUuPqcJuoad
ylVplwN/ca937XnVrjWJypliQZ4MdlJ7XSVMwErMqvKTQBy3C7NF9IDPiOtrhH2AAuu6UUddSgXo
OrFxqFw8sKts74gkHX+UgPFuUFyrbUxa/+hlsyDIqqNMbOxaIvt4PHzSe8LLD6g4pNhWop0yFcFe
YYf/pjiTOdc0G3BUFSDhPZlf5WbWgEw9aXMuuxtVa1sjIScg11HiTOuWIjkSgBM2qrz1sGlGiwdc
DrSi8aW33epE5GB1BPx6KHRYdoan6FXsQk9dW7zaEvSkts3F2dy8Xvl1sQofNrrC1EFxfzwN7gy7
45LlDnXLXLB2DI8KixBcl7OVW8ock6Kh0zZTkgJ9ZLhoD/14NcPCUX3PlEE1Givuxs7s4xCz/Y50
eVB2vINbeKnK9QzkH+HCyxeBDR2hfgMCt1y95/iOzcTeHv5nLmkppXV55Ctvca5DWk/DzZ6lc0Vn
osHdD++SHPW8hBnz5ahDH2ZVXAPiHgkil9tSF8OAhxV6wkUh4uqOZKQY5NKFkClw06PNa2jh89NE
UubB0ni2iLxd+a4FmfKJl/9FaHReAywMPydinaUCvnyhFgMatgsS/DkqXKRCV3fdlJBHdK9bWEy5
/kWZQeaL5EyMuj9oWLMuwa7EI/u+voJq26ppDygUnEDdvM3PLh8JcwWDDK7aJTmP3pubgXhNPKfj
e8CmhDbPP6FOzS/Rka9TQ+yYDgkwvE2T0ijFB7Xpd9gGXX56hijm3fydnv1Tu2mlgCfpZk52r6Qv
yvX6XztRy0Tmt3GK9sKPX4J/sdf+YGFAF1/v9f9Vq7x+dtxXuvJNy7GczaP4/13PJQmCFHxc4NAA
XQ8FRNYhYJNY2cSB7SDdwcewm4iHW0yh3i8/8Q2ENu9qwqOhfVRXOMnwdFX+04YaeQ/J3MNWSfvI
g5MqBjbtIVunHIvwRF/k64vmlixqZxv7C7sAaR/noiK1ENzuqe7uc7/sb4l7Lz7SkUDgmacnTd9S
IACIhxih82QsYg1v/nKGl6+3o+jKGP2Rh/oJ+2EU8esXPPL5uVVjBK41u+3vWP7ptPFvNxGJ3VAm
zqHve3ZPbS33UeowE/lGGyMN29uEOiCacMGB+99p4FqLvsIEqfZwjMM2nQrQbsgwiqh/7vDMjS1L
PK6Pd66XpM5aTvaVtaLe4nXIaDggCxpdCNzCm/MlgbiAkCReT8rbg2KZ5hxlA+yVZNHLGCdpzRus
Ut4hcYd/B60ZsCZgnWW7u1rbP4PV+2iEvaiylDnQykshMM+kFiMhT7xPy81KiIyG/zMX/T0jf0AL
mj5U5tpR2kiKjNg8nQ7H14o/buYQF2vqq0fkeuDS8waxSELJ9avTji4c2qfhSKdTKMmiWaTMq8a9
Bni6z5aMdDiSGs2s7viYxGGmoVcZvXWJcqAGNSnKa7teYtWksQmfFqdtssdm+MtJCDCgXSppgsGA
OS6t8L3+El7pi6o36YU4OcgETUdkQzOP8MSSfioRVWlNJcPQgnzImFzcUiSCRYVt10oYD3mtPuie
6LQl0Z8Rh5MjcwGyZ5iTh94Uni4EsOliHU1WrgpSRGrvT1MT7l2+7nGFNrQ9GnbWTmbQKawYlFT1
JfeAHSwUDDi22tMsNyUQYv5lOu8X02b9xRpMRre8yQiWn2IQUj57Zms0007tzPy1pK9GMsxb3ihU
5EhYHFo9BKnJfuQXIaWF16oMGIA6JV5+rW5dNk7ypwMn6uW6m1SKQTMnj12mAEPggaGFhN8aJ+Je
KjcG1CVIKbEDvuEn+b+bgjWRsW7DmlAEjxkCc6KHDodeCTb9wp6pU7xQeC3RcAkKfTeFwaFEYFMs
ECqZDqBsyYuQojx/hjnZBsi9GNaro9VC7AgqfqO7GA/btl44LwNVJQulyP07aDnRqzR0bNsmvNAu
n0c8ODUyK8RNg2MTSpy3HbI7TrG6Y1IUx52kGbK7CgKZkuL3/5GpX0iKVEB4lrjivadN87VAwm5u
Bl+2l0N5ngyuGfigSfiJhexMfJSR336YBqS4bi69Kl5pje/WgG6fzU9NpvFfKFVYfzI4hWe/pDly
IdVtzBOLJEVMT4DPWQ4fy0dlbHOUrsK0AGUzxyvKUdWPs8HahtJuUKuSQxGcMEu8DB01prP1KBAv
5sbx3sj2lDfcMkkourOgH2/MrjnYqHhX+nb+Q6y71jTFhwdpaq087YJkGi6iZ9S2WHh5ZYZnCKzN
PIsFYEPN8zsdGptzXYkEOnwVhFEGVVPlt/DQcF+e32WoUAghL7mO7QGxOAB1WURQMV+FxvGNCVOE
riTT1fDgrkxW/4noLZFbiu3Pt1AjYmD/JU7kF8h+rXZ65Fg1CMASjKH9GmT4JAJ6ADUUgBLiTXuj
3m49nA2asL2nQKHmfBgea4Z7+0vpS1gsApzVrCg1CZGOgx/wuFn/hjMC2KDN0AiMrPK/onRAfy7x
bdbnKyjb4sORNc+NvBgDh2zo0O/PSYDk90L6eZlTssdNhiW0bg5k98vAQk5kcn84Ggczhi3e/4zN
ajP5ONkeYD/c5gEkwOea3TycqSjndM1mW+ydudOnbtPKWF5Fs8gLTvodhP6LWlf3rDYLE/4FSYNd
m6SgfWQ=
`protect end_protected
