`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
anprbIjnuIHISvJF9xhIpyTU434rZQIyY2T7w0qBu1FONcj0qxv8JENCWOTPao3avP8JQ1q5vylC
mEdeZ/EG4A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mTtjyYnsIgiG8BnaS64lZwqfKm27U2+ehY1w1QU1TIFrzG2utR/aHJF2rTNpPer1ErENgxU0R6Mf
xhfEs/B6+SDFTKsYNFc9OuNFcoPO+AoJ/u14o/7w94fViqlIujQdf4uhJblcVaxAbC4zn9BuUbnn
GIjAVCpriijhvoXcGtA=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kMcwwHVrWUAmpHB1hZpQeFGL6IjSMFRsgM2wDpA9puCtIDbpB124SM8XSjCc4ISkPwi/q1n3DUtI
3ETjZ+HaResnf2JctlK7ypZ5iiUulZoYRZKu7ubcE7GJu1ahRaSjNU3UzSErmeqjq11/Lb5nwMul
7WW0psCEH5R1qyur18I=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IAbHNgay/GIWCDSyIwjkLkblwmHaElcvj/8LIsKN3QlsrIXRl0Uv2qUujaxWmhW3+qqHPxx4kIeT
p2uKX7CMP+ORhnlU8DOYUjRveYgVEqPP9GGcLOJI5VWBnnMfQ6Cj5bqLnab/WAkBrAA5LaZHgicS
qOmV9oP0LdZ+U1KOAD5/oaKm4GJg2AzO6D2R0cGvLOivImfaKJ2qCast9n4RF93Kv6IZY54435P9
Iws+xXLPS64Cvfs+tvZENs3dGFB8R/9+lbe+Kpi64O0fVAC3MvA3xkmr4/1m92qP48zzneCMDyB9
prjDVeqa7KqWaVLTOLcgEp01nzk4otvFjrW8FQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TkM9QxHaMk7oZ7fmjKuHhIsx6aah3bQeK/SlmmWQXua7DrtBRuI6aWwWC3wywM3QtLCu15IkMOre
f0fsVilApJXXbv0eoEwzPM2ho1gD/vUWhitPHQ/goIBvSe3J75o0Sxr8OLeEfstIBP+/vD3XS8LA
kOKcte7S1g3XImF3TAMCnKUDk+OPGNVsJg9Dtfy9QfdtNG+ZdcuNPmB/d/CxQ1uW/eDx9gvdMZbg
Y8DQQ6xiqf6Uiy/I0K1m00LYU2/cxqy4pMeqi0r9OSOW619PHsGQs7xYs4/VK9zga5w6tpZNq2Q0
kvJWaTbdqw5S6bw1mu2k8F2la0hGRimITQpDOQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TrmmHEVLCM39ek/cnDXVNuJnElQOMHF7eZzv+Sn4fqZoZqQRSSMBv3Bkn2TMrtm0af3RYw0xKFzt
3Ze2HbCp+fAWccGk/WbntQoSj3cNS7iGEIl2aCcs3bNYQACOY7vJSjAH/nd17lIdzbP3IfysC7pz
KT8PEJ4WlW9Y0KygDfCaibIVjJj5r+W0dRTf+q5tDt5OPX5C6rkJhZEAXyJLQ8N0g8/SZz2jHher
MxgHDeB4BMeKZWtfMok5dUMjODIKJPmRqBp32hYHe56yd44rZ9UcrxG1w8zoF0cquHWujXR/Mc9w
y17Y+8uRpzYlZ8T+ujwXf4UQ87ZfVUCa8KgIzA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10688)
`protect data_block
rYq6kq8GcWFlo6R34A0ZfAUbuQeVxP4Li9GWq0OTbvIUFqrNSajluO9hdDW6M/M6D0CF2Rd9EYQV
vjCsdnxiTRpUMfTXO9X14vGM7DE90Xmy8N0KjfN3kLXMNZBno7JMcAIWD8G9tKWVd0Hrqsj2r0AZ
eNWIhzrRhBptqpliKYmC/VQJz+ci/HG4Rg+z+VDsPpFiSzgaK1zxIVvalF8u+Bl31dLxLsLBOK6L
25hZN7aXNPcdhaWqKt9yKd53HXjSf6+sKBIk+xhQGLSU8/OXJ1LtoH/EgzlTThFcgI+bQUZduPPm
i3ZAgQ06cf+ZS76h8/WvIWThLggrS87LVHNofICLJMta8RZW8vYf06/W2W6fOPaM67kDmAhcCuhJ
YBwYdh1VjbiQGivdJQCNd/z5dGbzRJG8Qqs/du98OhhTbWKQSLgK9Fb58xFE2P7snAUQeWlNajnE
e361xT4qtysxN3YmJhR7GicHMny8wMCfSt81wODyQw5d405u8cOdLIvOgUzc6fphtVduFXTVjRT0
pAaw+6KvYe+yiRrDjCgGxu1N9vfWnctc0+ckFYDNfGMXlEynaUs8qAq3pSCIjeYF5r7MRZbMhZAg
5Joq5TnyIZN0K4hcVbLmeKzcII4vGog3lmXX1Ii3RBjfLvWz15cy3SnJ6marTWXik4D3lKdFRy5I
FyUDZnup9hJI+ze7aCAAkJZyQ2Qn7jj2mqDgysZjG7oMroX/JLZRprBy+orGJYcgwHxTql8kxLyu
UhP9niGW93r+gQBsyehDq8QKHcOGT65a+wrZstYxc/J3y8hVUCOeSlQLjV2EkR8oy3v5XwFRNPc/
aRoBLzKS8u5/Fgd2ZENPcCcvYP6Br795Xh1g5uif5dJwuTdDeZ2KOaBzuZaC6JXuLv6ToiPUUzg2
rwo6V/PazcZaO7MLH4BUKqABAIMvyN1ysbfp7weuz/Yol7W6fb5O/DXWgJQ2hdJXEduGrsSTciNf
LRc9unnoXkUGA8bl8Y0QCckP1dEoQ8ZirsHJ4MHh3PRVc9NHpbTC0VX4/0aDR+AZsjcnIOAffj/p
mt5KEv23fAEhSWbehwDfhXhSr2x/57Q7N/jsPWSCxSr2c63q6rVroY2hza2vUwsaoesHc3jP60fE
CqhonKfq2/cFt8aicMMoQkMb5XFF/kcr9BpqCRxD6htUmgTB4LmktLW25uAaruw9JI06kVN9HOqY
bfvAoYaJwznf/z3LCPppAhwXHeH6Yv4iDDZO9xotBv5ypEQuuRwI523nOexyq8TlFqRO0vG9m35x
XtlVDQxLS/FmWwtJL4B1lxW16FGWgqAwo5PFSzFPGFJACidrH2CYv6Se7Y7+0fAEIPtgDDgiYIv9
+dxaC3MYlO9KdoOB3IAGCXYZ/eT8fdzsySETTurL5t9+44c9MYg4KaYcjCIJ0aoAEIdBQfo2cKI0
8fnR34YLJsClCRvgkl50E5wEY2A1N+ozyXLjz8TjPlvg3Q/Kuv+nEIWsOB/4//IyXWmV7dSWOTIz
oU+5f8vu4nErr5pYkYpRGY94Oe9Cx1WiQjG+t7ejQZuU869Pjez0YXbtImqBp023V7RJUKh73DNj
VeYOvgVUQrT1tG0Ruw/GfSZ2d5vPbbm9lGJNL6wl1ZZPsGxlFtIPYpqWofTARJMSFPeSq9dCTXPZ
QxzetHEMB+oy+FaahVdcG747WZEDpNUuDVFVEn8cu45pUtSrinnhS85WfpfdEOXsb125qkPi9SWh
KMTISfTa8pfS/A5TOHk7YRongbRHDgdHvGeMBQTgutAvo6hkFmFB0NmwpWVUPaps9ujlem1z+pmQ
neBQfw2dLQzMgeCJII4dQg9rjHsccidcw8gdu3bHsYtmDN7Gqom+vP99m+cRTkl949lVdKH1/G5W
CsT/Oud2/oJg4rCPAABdHTPx6yovCY7pSwjcbfP6/PIjSoHY7upBcwkpVHUmchYEQtaUt2NCDUgk
J4hZdlSL9RBISyCpsLaYUEwK/3KkacRC3xBbalJl4mc5bKJrQRnNGTwnKLa4jFIcvFkQDEk1uz20
tXQGzXnvB/QexrhT5k94ernTmdzD7HMWl/HRmgtbklPltkQnHqC8Rzpf9uxOacKzwXP/lscPnfrd
7z84+z8hCkBfzrQWo0CH7+qiFMjgF+qNfa6Q+oCYS7wm6b5la2kZ9UfolKEAG6yNzrkV/n+GA/Hb
3GzwTolaesHi12TH/GQIJ8CDRdOKBw8XSIqwEB37BNS2gHyPazWwCMJG42uWnRuwQI5C9Lqo7lvD
0YySnXL9Y/sQu6JtzecnBJrmDK+yUYfBx/UinYzhaeFHvVOOeVvYFJW8dmCFUJQXWM+5PpeLQqfI
++UFfycF3/xrk+JB+xOHJdv0r8n6rb4Fu+vJBvmxMwuGXXl8AuurU960KZW1N7SWt65tNjvmNmqa
9MCiEm1G0lKQCbUFIphhlSfXJueDQX6v6o0Osb7t3sxsQ9FtyPBwqn7/xaRdpjeL6oyUKXyZfcLl
gllAxa+k/u4hyvRNyOuw89DzKbljWcW9NccSErftuCGsC6MhcMPMQRSpi0pJ9CbFHjHB54Bihki5
MscTJTfF/WevTmoItZSkfwb8fAFoIEMBkLTc9o+2d4dfRjPrMRxULk9hADGwGrkx0ZSB5stJp2dW
R84vsVi8z9Jp0lK2sGMECB+M9JewVCPu6ovOdIzFQicAMzT9w9JtvWKtoSodI1+jyXPB0pj5S8kp
OuXPEHWGebgVUxukhhXMR3tZFmYLwYMX6gehmPKYnVTKT/8YP602XS2PlYiqMxotNAgbHCz2AC+g
9XLXolnvNE4bz75pJLKGD/xRoZl9/8lenkTPxCNhS7YhMX7ZpD5y3HFOTk6P/dM7vPcQ1YtdV2WN
2A2cy4f8IIiyYzH+QsTW9JEdJz6xV3SywYXUWuylQUbzw6GmY76xes9/g2frjFmDNarOhtQgQnb0
AV01PGvbdFUEHTy6KpJ+g+ebKJyT8rFOkoBnWNYzdggjnp3ldZUaIE8FBOv1owGBXmsI7yohpmOA
UjOKLmP3+r1h1gV/WUusHFcj+fXGjwi4pNgXdK3m+XH4YtjoNuIVTEYSWHPf7Oo/hUHBuV37FqFN
n2yrzhicjVv2Wujw0u0vgoTawrO/C16QSaCWRDpmr3alnH+7rOZN1hcctOzKJUcp5lN4aJD5bx+h
iliEKjZJ5dHengZ7Xggy3Y4vQyzCDW0gNizqksRy0z5QAbsrArYlIJf0+zSHRiJenwzMZ2o/4m1e
yGT4NQoUUdPueUNJa1c2G2xsfjATrfhnuQ2Mty/lMj4rDPuc+cw7SSaycLBA389BO0SRrmjg9QQ2
ENpR1Lx3Ggq++LkEUJYjSyohWO2/fk572BqPFVskRczHBbVPDJpzmmWXklLxYrj/aH3W0SI5Hzz4
cLJFPSLb6KUXEVWy9/+HkiDYklImCuh4W2LLfrq5C4Jv1XPHOSEzK+G+hed1ZM7/tplpgHY+5uv9
lm/6WFlnKpwvFiIWqCkLt8GCwoKDgJ9BVG/mxbnK46tmOOnOPHx6UqVYy/+dC+6H3ZsaB44l0vN1
fCstFqPdutC0bl68Ey8Tdc1hoORCYXA3un/Klxdu20T7mnhmMG6SnhFSmp6iVM7mt13Oxq5Xss2o
ZSAMA2RSJOTGdIlZQYDDZU1S3x3Zv76BGUdxPH42Mf4XwcNwRrj1nSYZz1Mmp5yHgq9tYt9uI5TU
AS9jraqD8olNN2RYoSGUpXzLatoIUh20+LcIvABe/ZlmB5w2RUuBsO+JjXk5udOatKaqmg70Kk7s
bqTin/4s16i2MbCeeT05E4/VS+nXf8knVJrULR1RfNB13sWD8s8UiCYip+bUY6JpBCKsO0SPqVFy
7PD0a6/G9VL+qNq5akpCg2i3aWcmyishpMhXKciibklTPtymO450CReSZ5ki4OwAJmudHDubI2aF
SfgpHwlLbkf+sXbXDtOni1ydFUaalV7lhbWDyqFXrjaENCl1gf/uLMUL8w+B2fWrbIfmRs0nnisb
L4+gA1Fgn8Vi74mi8NudqOpT2r3CkqVskNMNjEw5mDnm5f9srzCryO0Ha0GLA59EzcQ1JCRLb3Pc
LKPJ4TtwxMPSHhHZKLzGnlLMljnpJjzrhwFGviZVX/LLRz9qF+rn30YudIZ+Y8jDskV8BYDTG6j6
UQNt7wAJmu+Ye7M1T0TXiHhZ2eYCmyfU8B/EgLguT6wFEGg4tg96qUbTb8j4IXfv6rfanzNTsUTg
6XimK1VxH43js6zMfcnJs4Uo+3R6+77F0mUXRSuyUtZGPXYh6zsciDpDjgt97UBF0P6V2nZ+ccoG
5Di4JZWjpRfOZV/RMpjNbxctyg/g2a46vVlpICIPgCd4Mr9AT9KYwYnYclQqkRgMPg3X2kjd6lav
8F7PLcSpollAnTHEZlJ+gdUdBJ7+ezlO43Yg9kDfVTc58XpQ/JThPNIYcPZAqea9+Lzf1Cgu9koV
deSibsVvGESxGfRmwQwTM1mxZubM7CoYbQpVgKV9owWXa+SHMMmGPLJNj+Zw0aZRm9QS+YL5gvhX
zcM4WHSmqV7FbVvuFybsgmOZ8A26Ng0xQ5iiWFP1VzYx0hWPnQaW+fKXyJXb1Mdc+EtvYOGgrzRi
bTLKXA78OY+kIfmmoKbUndQT3luHOgHD8BFEcdDFal0B7HXmDoU1QkK66czeiEvP8t9tSnh3Y43B
L4oQUmCtlEXNX2rRSXhkHy81EtjyeqHmmM2AELJ2GH6pF3MjrNpkCkvGlYTgOwbOR0kQRegKpCmv
xNXDaAjMV6VacUoIT5Jn2QhO95woI61NAWwN7Ap4RsSWCZ44F+NI244MQO6FOz7urSwKw6+UaJfZ
VeJQuk1TgR6iYky2Uv/YiQm1N2XSVRuHE1O+m+y8jQN338CXPFAawX0jlJNzYLA2Coy5VZNiNYYh
wZYy0FIDdPtP/MT31BTvQOWQhP6AaTKfvHdHkxL2BGIecZcQmN69BB+SbitxvTmby0p6pbubJr2X
FuzAFfFziMgGg0Sj7SnIL++QpbrQfyox8pq0SCL3VK+52ZdDLVJju1EhR6jTOCEvvHtmZ1d/7+to
HzkVJp92kFaEN8y9AB/wa8AI4f8HIcDZYZHGAFldjW4wlpryrVQW/TUNcttCxSEbtTaEQoXXGbUA
ryiMub6knQimm6JqXrUt9O+ttwMMC2HjkRcYqFo6xm9qaKkuCXxAX4cSHOl2usBomYZdFpi9gXwe
kUPMwrM3gdj1cELNzUSf4PpuWcrQCUh1URIQzkEKP4h1nhHThq7KKE/xcJ6u6xmZe98UI/jcjohW
aqzZl2TW4Iodnn9ZKI06ZXvBGC3N7KT05Eq/kfbLzVDxhvtDrTjfeg1d+t99t9I+cOBP2otB+vze
hz4TTlJ5fNZdWU1gnRDaVrheOQF27g0la3/bdI281btu/gyes3JSWtLh+/aY/EuMYM0gUCadbxGo
KDIGG72cq9SGF6uAej95a3NRHa83J6GSeIMxsgZ8n5zYpLV/geUvNSA1srcSJAcTen4xJHnuI8IB
tALXZ84nin6ABhMmK+EUDwGNS7q+TAOkZyqi398lzgJ10/IZcU2gSNwUi3R1hgAM+LOCeZ2TeSox
UUPPYp1vjhBIeuST/miKrGTAzZEws05MDgAvczY4Tk4Aga1Qg2PfGQrfR7Rz0YndJJQMAs9kTOU0
BnRDiynpnrr3IqOhDgM78FEvRVj/nYmYXIm6kfNe5FCM0F4YGZ0HEgahMnzDmxti+XFza3XX8Lao
eUiLyGkXXSWjgT93mN7MKIa4jpxZSvThz2BUWx9ae3HcV2qNpMOGSpKE8CbRp/VreDDmrHb4cy9T
bCzg0ZdTgl2hvkoUigL4ETqBjNMy6XInHpsUmRN7/Gt8185T8zeIzK1kghRK64NyhqH2jAVe4USD
1KiNMp0ieus3bkl0IkDFnfPutwyWGnP2BVMZDF3NJvy66tCsT7C6JTBhlor8t7vb8uoqQDD7KXL5
x7wY+NLKA9w7DcXGey4YPCmc79v1nh1NzZBtwl++QSEA9941F7EWOMRbvYZqRGPjRT3qP6uDfOqg
bbkaooZbQcvf4tA7jOROdAXcY6lXToUNyi2/fg0ws2bvZ6EggWWtmsRpbqTWExSfmIYVv5xGEVAB
mNORE5ziuhDU2M1S6UTiUNItCzxG6ws86ur6q4wCZg1sb96cO8fJJdQdPhGboUBXtbF+HZ72rL/t
5siSGPvT3MfeHzH898xLeqaOwxWCnPH8X6PXA2vlYEQKdFCX5kudK9HYa3DYGnEof+u2V/4cstLq
gwPefh2z5BG0r7uaVAFdk67WhDatc7ZLPhA6aMta7h8bv03KL4T6OhuxnxzDb2TgQYHDfe4lQhmM
aOJsywmYAGycU0I0HqnEkIpYgo7g5B8mcHp4AHgIvj8cYIi84ZySx+VEsLIBrsg/kVRik53YgviA
QoE5zl+RbQ4plJ3cu5pd9Bv7P79dc8ifcsOKSA6Pw5XXib+H085x1xNAXPzGaEVdQ613kS5dSXw8
tdyenIQLfYgoy/ZG6DEeB1sFW3WNAvu6KzQlt8MZXlYTwkcuxnm+CFdH16rYIIwjsCkf4QIwhAgJ
66TRorlXO7rZhHhlts0X1ciaNd8xWHkgJNpIrTBW7QXFDwldcMVxGOMO1TSEOAKl5QY9sT0UGVVM
6J6Tb/rfUg25mZvUwfEhIErJC9u3EIhLmaud5LXtEs5Kv1yimaEl/z4aD0+lGSZXHKGoVoWH2iar
zxqpKZB/Zc+TcChsUQdU0vYA0uldiY6xOl//EBZT7e9RA/W4a/98Vd8/OiwSO3XdwOG3IbwK8S9X
3sq5ODQOO9Tn2r1mtkVSk2glUHnZpcodbH76AUOeEv0W5tuMgS70T09kybx6IQS1oli+Yq6LcA07
9HJQiExcLxWU29+Vnj8HBPTpxlm6VpDWvu5bHn9xA8H9xIj3qVMUbf8WPWta1Xi58ml7GJewMnzd
WbXctc4dQYTS2Uc3ypH85owBlu9gyx3+AtuoeJzrmycxv9xcM+RX0fX2q3GtKQSf2qQu6qk3bIAX
tIS+kYt6SLGNEgSmIVil2340y7oBZmf+zURmPF1NLvNcwBVHbK3VMrF28OrhgfKVq6GpuqAiLHcS
9jQbrzLWzqP6fnBBa2d6cqntJjCJmD6g4rfZIJF5onIClz3wLV0HEEjfAs5j9LgpTKfz5eNOn3f5
mfWgzZKBtj0FmOp26qhdes8nCzXrinTFLRLo7VvGOiorV5M5d7r+Pw4+y/i/uqJziysJ32pOFrue
lsiBgkouc4vz5BPBdFcwn0rNrOilV7gMje2toCWgXacn8yBM3V/iQumuT3g39yClaKsJ0GNTs6m7
QPbLIFKmPzIPy/9pJ4sIVdEupg4KUhekuiIbyLVIOyftKJt13TJhtDdU2TsZ8Oe+GO+GRjvOU5zp
44A+5Ab7t63oJxSd8+9e95wYuX+F9S25Q/+nE7B9CqZUJEzTEEEdpREn8w1AnUaFUMVzdZHquuDC
8n6Xwim0PcLgRC+Z8wevq9E6iEkiyWxLrGMUdo2aP6N3NEWA+xQ+S9zVrvEJoii/aNa7XjRDTu63
wTtD7cKBaAHZJQlT5RVBm+tmFrxxWK7FAfP8eXf5F0X24mOZh59DVHUmIwRP/UjFTuQmJ2uUCqwT
L+e0YQrAVNRT4j8wdIGVt4rfOzHF7vvMu75OjnwT3drhAMtBKyNBb+GPdy/UXNf19YSQm6+MH4SW
9sTfOSJJj+fNZzmzeIKWDEoa73jnl2vNfcLp7+uX48PGmBU0U18Y9dYGu6jFLka9Skh3bL5u7+VP
YjxFipcFniLlHTgkBSdKrzPsr4p56MuCW87kFtItW7v4a+YqITeBklhyFEwewE9vdBwwO41FqiBV
XmT6fllTRRW1xIxVa8vV/4OtSlfi4ePt4cJogOojAMBb4jzGi4451kPhV63bE3dz9imzty114Ujr
jFsL/VF2sJyWo6zzbxyh+7ApMHEo/EMGiWPGmTKmvP/XbasTts0QqSDrjvo9K9qJx8S6edAHkxl7
Oy5B90bWEENdxylIy9NcyDGv9j2E4R2OPHA+jlgXTLJHP85Sk73SdVuRl5vtKQZYxaLQXWDzEAY7
a+ouo7HdeljiZumJhll17BOl5jpp2yPN0mLnZABU0rphpXXIkWBXiZeAkkUXni179osQHYNreAip
KQV1ArLG6K1CGxpIPJym/FxGCHUQD5qcYGQIa+25NIHbAHx3pDROwRt79/o1SIqzdXq88dMGpSUi
ySDJnNyphIQAuq2q8juegaqrVoVKwR42wkoiAKKHGqMxRLVeL4Gy/UUBbzrWPp9wXGrMvy2KkLq3
1hnUKMhWpa9qoQ/1f346nFJVFsHXeF8PNmDuEHC/2iTBQMvZkf/u0AxfINVXGSJXNmu7AuCAZN4C
vgd2ccF6+BZHrmsLrZvClsowoCuJM0CY48Jg7RDflJ406ETG43v6eL3j0XU7I5Opv+JGFb5UF29W
8JWSjIA0LY0a26rAbMqYoPDXEcOVdRiQui0gCvMwFPcKLtUZJg/XLhFBw4b2TX2hY+80U4YexF7G
x/Dusw0P0JkevYYnUjkN7rJfY4BFbrEhxEiq8DOYe4MNnNNDnqZ5PnGKMLDwEJRTvoTw1k35ukGU
u14lzu9t5Nm2HRZli2wArWmYc9UUD8C2+zoro+NluOZyTgt3p+WwbYxr1CoLzxyKdxcFZo2i9noW
0JRB7Q/gsTXuyD7zmsMP02Wm7LykQ3Y8EabAxgXTS6XlO0g1mKKSIcVd0IueauHFUaJSP9XJZP8o
lkNh64yeTUhEMRxq4AoF5J2FH07jmbHiM1DH/v/G8PH2aD7zrLxIGOpVaPArCR4bWSiPnXhLJEI9
N5OtFl2kDuj7K1+9+mHcc/bl3ZNyN1TJxQ7I+/YQG7EKzDMDiz8LlD8SOP4nw/zNs8Kw2+whhPhU
58oh7SAL1g7kSoLDCzv/4Z75qBUcG/WeL7js+y6zsS7rzB4DbrIq5TLLAMzVEmXjK1VuS+Ttp4JU
Hu9G2ojxr8qsk0z5wJsSw27tZkaZ0SraqxW1Qq1jmwZtwzi9BM1/GowG5vKnTt5Ab6cYLyzga1rw
bL0/YU733wMwu+s8twfwhePXuo6b1ZYUJIFaxxRbmkZDiHhE5RrBio/YBVCMfPsi0pKH2ZCAFRs2
pZh4nSo1OgC7GTOYT14V19rFvnz/XlGmm2sUG7zCC+uwFrbM8W4uFhPF5Z3UspiifOHmdAl3knLe
qsqF872qIv6oKaO1Qmt0nwVITrzKqFQys+9x7aB56cvCg3WlpR/vsoALZXSx2nYDVfuJUbe8lnqg
QSL6asb+Y++zwv4TCIe2UXTsn6VfT2afQ2wmmMnyxCfMUxD/84cIxg33OPU3oyuwQ+JHwlZ8ZARC
wC+1hWdqVW0V1ZJ5m8GsZzBm56tJMiXgOJv+cNxsQJsHsIr9ppM6XJtkQQMqtb3REyhGdmQCn442
ARQ+KXsMT0vJHJ1/tCQF8g6k2Wqkc9zYK0dQdKZe31a0sxo9pSth1gZEr1YwFfyTD0uXxW0GVqJh
8R8z26RfX0oM1sDX9R6YjJcaHh5ZEoycQBYGCHXs8bLyDhmSnWGxwkMDNXTC0ywx/ObNAq+0iTj4
KikdMQrGYacRzmmAz/MuLoWynkhOmdg+9Kbk3kEbPD3McOy5iepJkgG2QtGVKZgZWw7gSviP4f/h
1UXyHyn6BaN3VRfMUtMV5RiokWfAUU7KmsQ2YO8vuLSOUI46q0zwdELmVAAch/Zos3DFgysYGkto
vu+MvGhZJ5leAhF0IY9vMeL2GI09Gb0l/3AOUhFvzZfknjfHDJDLwesShKWEikf6z+DRDgtTd6Bj
P+wdMJ+FZYSH5HS6G0pNx2/j8ryqFimtRzScfrGWr0+xjr+01MDvej9PdtUD0vQqlaG7MLwIV54+
LHzgEUQH6ps+RjkyZgEFxWdBuN4qzyHma0GR116NxTJRwM0ME+yWFEghz5i0jsCrQ2AeiKp2FCKk
OWhVk8WsXxffYllUyWw8G8xqSy1iPJegcsH4EbPozq3g83h4Q+hK7uRvmnZiDCCSeg0iitrBd7/P
5LsmHfhh7mYLQRVw8nA6RzxmsJbEhGsOdh71ZaDvOYaUZJWCm2zWhBNS45ZcvrbD6+p29ityWFL9
2Wg4GMr7I+eByaXn5+RCfojD+VUEdERIuXXnumX0yEBRyoQFRCr6w1qhvk+mZp0eefIzG5d/tS5Q
WYcowMMjCSbZKmn4/k7TvN5QTw6OSUGrt/24m2KSjLRd9gyp+nVAnIPfNlY+TdvlaYYmPatp0F++
ArQ7I8PhdEZJHsd3fGjbXaBlRpwoJecdIGF8IiaPNa9j3n/ITw6ARxmPWm95uc1I8uAjVDQYHTvs
bDw8SRsbHHamfdIws1WQqoGvm47vejqZhvPCTpQ5kAvlLRrcfMKfm8bCKJjp6n/tN8yCfK/BfdcE
jxBhpM0zKIZR8ARZ1kARL08wCga/aiFi1XVaIYlxM3QIVME/nUdhjPe0jafErCfhoOymlgWc8hgk
G273NauBgQtvq6fkUZPrN1Sx2AuAP5nxFc2MDykhxeG/CsZihyZU+3YWz2EQ7yd4xebaIWIPbJpw
zAmM7RgE7pAdW7Qbk64xb7OpHGwhjd8JX+ApdHavum3jVbz8fDnjffXEFptktHV6qjRn4e7oi+yo
x8R45J6ZNYhigRB27ahg6vW9JOH5yXSNHpazKX9+KWKxxj8WfWOUFEDjsJzlg/nRjz9blObC2/Uw
kfRuvmeQFMCta0OMVSgqvjMwlTpRvM4htOCkUVMZpXimPp87Sk/6E3IKyB8vaD6ZbXdOAgKuwMmR
eVzEa5cOfZn1mztij1XvT7V3pK1n77+TihSkgD4V6AUT+bGSUk4YV1NYHq6Guv1NsTBcS1g3OZfl
mTit2yxTqtaQpZGk5b9lnrnx4h9qu+vtQA1Nojq5s/3W5CgCjAJZMGtuRZEpKKHbVqU22DVuEm5A
kltZfn6wmbBYdwSHo2OYLxGVD54Wk/825MIbtV0ALUnz0eQYCcCIWcevu2Dwrhltw+ZvvT8e1hAp
04hhGTwg9F3LjDx2iuE7MXwcKaDf/SmjMmJC5uI12mSytBSQ61hXrFsgcnIEfCQCMBZUOB3a78Hz
eYbetpT8QdvwzoXCtf52RH841yHOcdHqI1tLlhUUxSIZr5Eu5imda0luikPyUKONIaf52pCl25Hl
LDtuZesEEldT+ahkFhh+wqtAmYLE4xycSprxlcTE/pCj4FBujbXe2gmeq8z+/A+eP+TgJTtN9uwg
g86PwH2/N2Yac+mZJz4+D3C1fi5pVhwtk5nXzaNmCjaUyJiUFtz6sng/Yx+hZ9qncMAsv4kDQNIl
/KXyPwVinQzyq5KvJ8xkg8afeb0J0JERwkTRBzRsuourQjmqF/AqUKDaSdxf1JgT3b/gdkLnaLtx
CNfbaC27kF6Htllg9dVdH9LwjAiI1OPxXNCsbl+fGeS01Qo0/7kRcCFjNXHLuDgzRvgD5gJsGWB6
mFXkCdYtCjlHBb2TjPJFmRU2mM6UpMycMt0xhuK1CZyjJjSv1WQ9G6l5flrgW0HxaqbjRLtH4jdx
hFb1kkYqIfDuC+4p66Q734tId75Y/0TFAqTP1Uni3bZzr0DZF+M8QnTyystZjQd26jw46t3yc1GO
Ew5e1kt5/WyBkFcX0GStoyggflpfvqekkhhHyasGZZ373f4sc9cUq0nNsBWcRxNkJD0pk3VbWxuo
7n2Jtr3tUOTCIK3te/gn9553WgBRrAUb2x5+oGNH9ExQwtVvpeZzHLkH5Yj7VvH5aV/FGjhExklI
bv+JATX8XG/CPvYr6/p5Smi1W09H2+B4SD633jpuzDAIRN/K/G1jovqrQW5/+JOpMZznVgUaf3Kh
qlMySIhP/J822/qc9RgjDIAE9XXFeeNu9KA9WmetbAj6lN26Z6GUfttGpjtSutNwjsBBsWtAFfbS
0uPietlNxjMACEeQLiIf+Fb5Z30yfDpFN5qHy7R0GMC4Lxh2HQhjg2PRkNXTas6XeDpqb9Rpb921
9uGA9Nm+71r6bqPs/3mOcbcAWqJMLBAAVm1o19Ea1i8QVN3BGqKuv1fxdGJvhnotxVVauuiellTt
4viaPsaGMeQhXgJUiCIP7njVZNLbba6v9w7fGDq1R3kFOh7QkZT3SHU9AEQzjmDx3rchV/1FRUUW
U/7HoeUlstoxkrAtZq7HNq9Jw3hLKRAuJTW6xVIt/geJw78TNr7hNCuDx/t120FxlPDy8NPBCo6b
PokrkRbKqk4KWaXmfNg8ZhgdWP1xRGz6bGmpHIjnlu/dmM5x9sPwyRQoZ8jatWBasBAY+0TrPhbE
h+D7hg2OeVl6YORWPaYsM2w5oDkS/QEcc4YVWQ7s1CHyni8CxRhV5XmuN1E9pnYdO6EKEtd0uJQs
jk3nFDcqmJ6Cuv4moSOXFyaJ+fbTkMJPo50ZjuN38MIUk7t2Aat89rGFRm++R1g774rH/7tLIjZ3
CDNXJIjd4kqFLfSydB/5iZCBexGny1jbWspeuYBZqJFcwVdWo78kbQTbkgGPS/+52ZLeO3CAYd0e
MTYa1e6QRrFQ5dSvjA2pvByZGHh9jgxfUgOZk4m5Zb5Z2ljoV8/7iJ8rNYzedAnXB5XMciwUBb6B
Ue/oV+MxeE0U9XopVtXlNifkO5Pe2ioT2Eqs0m2WKCMUIznbhlMvMRdMfqYs4/dg4fi5W4vJ739k
TnbiJWMJGPk9D0o73tzQxZrAsruLgYy7jLjV+D4TvG2+p2fkqOShXFF89K4hJr0QBrBBu5P/9DSZ
JAmFP0VkYcHoN6MN47lpl6nxUl8mkxCqcApsvbVkOIHjkpAo7UE7uwibnXjq5WGGom4SmSO1j52d
JzJ5KUtekwxNaPnYN/3mLuNURWnIwa0D4sgiabLBmfpRlC+D2G30LMhUA87l978viD4RRZEHKiSn
zpJSrRvmk55coRGi7uYTBtAt3KdnuwPmAuylcUQgJP2HMxuIfq6GmYj9JiHKCa3YwX/piMHAu3/h
Bq2K/wbfpf5bkEX+Y53HVuZHDQu860stwBUsodN9NjxehXbbxeQXRqwTrtdNtxb6+sBOVvCB96lI
sW9lzldswBnaeqCJRJFWXR9pfMYCvLffFAR3Yz9oFZP87SBScWDSJQeFpaurtoF0LWLIhwjdgYPD
TqYtDYMbPG/OFibMM8TkrB910APa3fcA71zxF7qKaIcMfbIwucGKNuaAXg8xL6cdCGYlJsT/Mc/A
P5g/BPqtJqI4W3TYRXL7Lt28qxHaWw5Mo+AsIKV5EV/s/i6TiDAGiGC2YkcEOwF8QfJ4HtyaNiWe
kiExQM2vR8+iL4h0OtgotVqFNOOVbcy+R9sg4sIcFhjbXqckEE4D5ITaaJ/11/6D2hqqBpQrh9mn
QXReL7cEDUgTrYKYOZ9kswhdbOUHG/9UCLq9z/4oiI3X55GF6wgoxhEM4g7nipsXEmzAjJ7x6844
PCjgz9cAiDDyoXZ5bX0mHiE0FStgwDpePIQCuPbdfVKbd+q6Z6bEi9r4mt/JY91nQebnAePy0HTf
IlbVjbvC0slo8f9IZqRPt33z0fUbZhi5LjkoDwyW2QWKZYPJNTzrpzrUvZwwMbbLvn0arwhVZmuk
eUc73yJLwd3Dund2LjzPGBaXRD8xXKSOEL2pQcYGfyTY1F+w2DpwsYXkFojvsKt/+aRcwXUCfR9T
YEjmbhTd/rxLjM93fPUiohaGRkE8PJ6bzqwlT9b6+W0ES+GLrvRpEGETDfs0GDcVW5v1f77o+CRd
NzTib1nofP44J+8OSpyiNGSEDZsobEmVJ5ieZ4UWqqhKfwVndCbxnKF8CcRlhc3VdvUNNOne1LU0
Dn+DfUDRPFqV3lZGn3rHCmfk9oxSFfBGhvSJYMIaTBwzDSVxO44vtB81EY5AxGpzJ1NraGEl91oP
C5FmBABOwPSmT0xZocrhy1Z6/0dlobrRmHEpOb4+tztPJWVUVQkIw9VnLS/j4IoyykncD/H5G0Wa
hg1ajrS/PVgo9HyJXu+OaBYzqbmqpqBmX08Xdv+2Ebd37xZvkN7TS/yM31sgWi8cpvxE2PUXY1iQ
yHjALphAtzJPlpgvWn/WEulboYY75BOjbRXAiEcOCEoHkwahvGBmlX63Ac2yqPKWHxgaRPdyjI9x
Lo7Id2z6UczQ0RegLPfmZoDVToMQTmxpQXb2KsM=
`protect end_protected
