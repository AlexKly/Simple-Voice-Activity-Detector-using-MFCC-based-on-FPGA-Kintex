`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rL7N9PUVRqNu4FFbRGrHPCfPH25d02HIQlr8y0sZoNIRNsRHLwJOWPhmp06T+FQ9nieZUez9c0DB
8UfCC1rj5Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KZcTdSyf6a7ypP37lt8e7JitEDra4QQQRt5ls6cgix3pMhdo1DqVT3onwqTBtFZ3KvE5O0UeM4x2
fZHdy8ovPjQ1uNRUwZ0UtMZdJKNzqZj8yI4Y3NuycoU0a5A3YwMtupxx5N0DRzWHY/SuKYKPcIzz
LL4a7rmNXh6vuNbUyVk=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VBZ18aL1lXX83ZKZMPXNkaQCX/HjjTcHVdulcrXjGCisttzzLrsrk0V2O/gItLyk84Ql8LsvD2Eb
A2O8cckJqLdkHuaxltDeqE/1CIPYed5QVIrWC6wV232PgIpW65ONHNu9m4weoJ8i0+ovSid/wNpu
fiT/efY+P/axtyDCQ20=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XBH79GRs9hEVvuJ8ooPkUcQRons9NJ1Yv18XcgEfKj/TKTvJtvscPO/+Nnr1WN7+HczJmkGjDbVH
Pe+sqGAyOvryn9uJodO/TT47PEZKPg/RfoD6IZIJw/AltKwtdvtHZwDoB7uybcwW0YdzZLCO2Aev
fc/hQdeKLPUT7qYkUvGwecvd1yA7JYA/NrWdgJ4oNyf3Pzu8dS/O0hkazYUNNcTCs7DpNF996/Fq
48eaEHLN/7AlS1n5HCOVknBJ2GDD7Xo+nI4EBz5lFxa3p1kd/TDW/Jr7mZB3UAiGtb5IvNscGpFO
ZfQzasfV2pCjXoytQ2oz0I1lPYcQ3Yyo7GU4FQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MpD7YP6FeOHJSI6xynL/SjzZVdA5X8I0l2D1UxjxWfdBEyHYPHgpkgY0glHnmzYsPFc6dg1sKusL
vM5vu45AoMJtDCKXZzDb3gDh4OA/A/kAf9r2VWD7HnMUG3RFn6b+stlrIWiLeVFNcbu2afHptHAR
T/t2RivsJse/ls+/XVHJdtsA1Cx+6C11KJeIjxuOy1v9b8JZ0CVzmQ8IplY4kMgaKGkfu63+qDYq
tQYqcIFyonR1aCG13Jc1rxq7x9ni7iWefWN3WjhhdpjqJj10qgv4Nz3Tc4YqnmOjAOAYODolKd0i
e2IvYqJ2bGiDWvRGbCxuKxL+7tlzBkLiaG+u4g==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XBA6eJpnTU7qcMRnCubuHIqSvD70Z/pBbP9x7EKiDrvtiD0XNx5yPpn75PzN+69aZtGUz7mBIwRu
4d/QypJfep/6rPOu5uhMHG+ufv3rhPm9LdbcvLAKOHj8EpkmLuptLXTAOPJjlBgG1V31Vymdtr0i
3IhyVOXrdTNBu6SmrIlu7hv4AII3j1cbCBq0cKBrpitPG3G/mARZWBMs1e9cdgsHngTd/XHOPFVA
ID7ZirMNl0FotJBylf63TYsbwV2tYUDECvD+eD2qyu7U8BMZrawKjsy1iR8lnVcrJ5sgeVrzpkaV
WJf4CSFf5QbCCxdfuqARqCp14ULHFlY949498Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13840)
`protect data_block
OkuQo08roiHgdZG8RAepEZj65F37liVVPoLmqMLPEnXwh1dd7N9eznDXnG7rUDmeqWlyybdFpCVy
6ghz8XQTxIrkrpKPuzdTmRD4iJK6ahXaop1qrZUfJ9GU7sS07cS8kNfY71DD4BMQo+LJcnR+Utgw
PLsRO8OAAAqnUqRs1XYCiiPoLtKLbI22FDfZoKarniN49DZ/5Yj1fyhLBkCFcrA/K0990NWmQXH8
J/3vn1Tv3PoDWa4JgMOhBiLlqK7jDuol8VZNZckijXAeFmQ1q4VCUioZPkZaoZdzZV1Y9MbB9IVv
56mCQ5MkpC/uAxYAohZHFnNZnOCJpjK4PanaiBpeKhuToHzaidGlySsiiTa9KKBl0D52hoWvFDSK
H16wkCrNk8T+GE7oDyTqGrd6tljHGfjGcUfysYt7Nx3dObPX454z2KPEWd6rzM2nWPf8iMy+N3dX
wMChdm9I6SfUoPMfgVYdQOC46KIVH+aFMa0G/t8CllSvWxhcyBOI4ihktzlVZadeIp5esuVYmvt6
tqEGM88+oz+yfG1yt9Vi/xre8LYqa0jD+kuYyowabTvjpPkmn7fd9DnQvOJijG1v1vOtDJcleJn1
CYZrAzeIDXme7vX7w/WfAzLNYRvTo1cWEr0hhSURQoc73owtC4a2ebHyBQoZ82jlUUXEU6TeSfWl
WZKdjbXuy2kn2DSZNVpiDsXnPcgbmvJlNPXYZwAaTfTyOY1nBE8CxhQ/4ThzHAniEipqzdAjmyyj
3AG91Cq7oX07/h2FALccOGsU2D8u/ZquEGROQ7s66FnJH4pf0Fy8QkUUVolDFBMvVlbkRqYpPse8
j10aSrjPJa+bxv/CyuAf4vV0N2NX15IlICQ7tOQjFzhxmuIqpRdmbMfI4ahXUNKd5OJ969ZJfZjM
VpHGExISFV90jSV2K3qSYUNFSsihZUENDXWG4nz6movoWR7oxQhplykHy+cZMKQF1uTQzUMZLfQD
El3Rr2wZprK2DrGbMuR4XB5Nad3J3WQujBfxvS8TkYegHL9ryUaiEo9J/xthfiweBKjaq6DA9Hc1
ipvViz0h/gXRWpt3plIMFdK7tqYZvu4X5TOf4ufEW19dqfiOnBGpGdOY2F/zv+esPDSFVlSuJV+B
yPR/dAYI25WYtxM2197wPdGpfPBn6EyvPq1V+NC8SVbvj3e2FEQotuyNMT2dnUiKssNHZRvCvAxa
Np9h+/8gbg0crP4BMNRCryB1BvPe6w3pUmlvwGXCLv41c2z8vAYhDv5CH/kwAS2JtxQ9PlrgzRVb
13LdKdrbImlQ+x0RtEeDehmq2lJY0sqBPvratgT31p+aSvjUNiV2yaHNUAugBOqk+g+uaCuV5JtS
uO4zWlxmNAvF/lfVzcm6Fe/LQ/+SnAsNvFYzGy5NlsCJAPoh6jhgObPHfrrhMLLzJYcyyfnyXc+d
7efWFUvhan4t1rQDDBrpMGHc3amWHfjUpiYWeitursB6ewD96gPlNk9F54lG9lIaFKLLts3AopNL
b9i2CZQNQc4IXHox12fXi3nASGt559pzcFQFiKnJL8WFsOzWLXLHq+3CHkPw9i/HCYqC+O/lnEo1
J5FGni+R5JB63AWYoSIqgkWjdcu8QhIfFBr9JAoEZD4Qo1+t/dsy8h3qtY19QdZRDIf6bykNG7bE
4YVKEc443h5YmFbaYSUgne3W/oD7meM75nTE5Cj6Qqlw3O5kwW4i+UGxPWUJxfFb8PsT1dV6iwj7
/qLPiUzUAKbr9um6oG5oi/VqzHlkGLQ1+oWDPPsqELw6wmcDFHfprCpkxdH9JIZK7BdvuWOR9Hcs
ayZxYeCD2qXYvj073wm4O2AGRpCZHFn7wUaHATHGVo+0s7GgVn91ymeHwisezztj0fWkYSqJzZ6d
f4uGkkn1mLfQDmoyI+tfg9Uk0R294FRIyL3vcnXqZCAD9lT2uMvppl0dYtmem8L5S68uXQzS14sQ
l+FZUvQ9E4ZKluUdmLEvcNGUfogxKZ2lMxPS53+94AUhVgZOx/eLAZ5OMH7JfuEPV5+cib5ubf04
T5aFkt8F5wcF+YnvqPkRObdt42WuuYt8bLay7C4pTUZSDlgfIxf93ketfpmi1+9EzrQ5wYjxtxDC
i/tLNObaY9Ow0XLD1H5agavw4VDYiniJlW6fQRYtCtVO4J1uF10tur0vrb4Xm3LvCqkcvmHEV+/A
zWL/o/7bUWVdVIiHHWc15Vi9u04WkvSXv0tTgyRMSyCAMLHVIaDUpo0sPcTpWa+UtyhUHHTfg6pU
VzBnSOSsl//vfby3VuuhdfpzXiZdStfSHcZIAS2vtgWr78pKksvbveMwpiaHFy5ghJO/xnmSNaXo
WmzNwZaJ+0iJeGCjo4IAMb3RpSkmpdLcTnGJLaLDNlD3W3HcpHo+P+yDvZKLn4fbqFiW9h9W/mb7
t66JPfGb/4EhmZLq8Bb+wjFWqcnHEenIhZ77SybzkA2UHE+B4/Qmi4Fy2oqvmdgh6KsV4IhE5A/F
BUcjJ6CyFx2o69spbMqAdkxeYwn1U94L52K7Ap76P9NWHyes7PNFT1i19yVcrm1PST2Y7IHj2nBh
NiVWyDFtoqz0CRiCwJkRBKAm8uVJsNu5wWG3O+H/BewJOGjqZhELbScV7+pFx+Ls0/xD5nR1vfD9
gz02FAf4n/hFf17234Xta8OUobCLlHY4SGTU6S4SKEuBljxejPcVut2mcDz2I1N3HzhVNsF1s/Uz
d7V3HZ07wvqUbgU0SR2ApvM00rBgrsz5oBkl9Q4oS8j7exhVqCxIXMHXVRTh/9mcVw0ITVk4W0JG
htrrl2wWJ39cvS0AWdKMwmYY/pljy2POACaaOUyYj483miX64fzGYO0bTYbG1PWtc6ed4R6ajfjO
BhVCeYHQBOmmqbLUsnrKjT50dALVwA0zGAO6oDE6/ZKkuKA+Cf8V1+mSMCJJ7NT7F4WYBej85EGJ
7s/6SIkhcilKNuKQYbP/buDVy92RmIJOUCYRujouyXmjIlUL8YKa3cWkM/2cevblby0WzIh2YmhG
uHdEEbpV3zNhbxo4W86LMuQyNBRPWZp0FIQQ/WTv5EiKGlgvRdK1T/R2ijpQv4DW2NflEuSxBPcw
jxXAaEsIRDbsTTWd8WKiLMLcRK8f7JaDSqQpWLT8Wp4JhJ6/gonXcLmY4bLxLsy0zVtLbbEDEn4j
6lFE3DsAY2kQ2h/4mioBok3CPMmkee1lkcQ+hDYchr84Le+WlqBsZNbgjHCL/UjLhhDdhxShe6f1
+2k+CR2tGAgqib8sFtadz5OoxZhwyM9zwZ3EJEr2OtKnF6DKVArKoF/WNCxEEdq8AbeIbbOxlu0o
rKkjI44NgOacNL1JmCOVLRoBjbH24ru9i/42n+LDXcWHyKe+NZEDGrFYBI+BgXb1gBQ0aHat+gj8
LWO66kbcWvcEwlZK6RlyAquTF/C1lu2hk3lXwXYjbLTFybGs08r5c8CT8LUglPTfbfCDnl6FaS3q
KvyxenUKCFEZ3nLu7oDD4NzN/dmPX5mgWx+HItFNPApIX9ZQf1Uc5Cq1zX8NQpsw2B8yo50VuOZ8
f5XyWG9iT0ru9AWcFmhhgfmHdB33aV8Ti2Vht3igCl4XOshG6Wq5EHFL0+zDLiGjw9Cqx5OVrNEa
b41YFQKBbkMaPW3w6MAD+1H8qylBX2ZM3RNBRpO3T17IrA6Pd9ITCvdu0Ax0w3RgrmUa1EUzHACY
NPN/57X1omfRztm7UsATn34X+GDHVMYIq9wd1v/8PpyEtm9T/HKYq/JuCXKkzqUtJmiELBRhQBgb
s9f8y466OSnZDtaaf53wzlYWTkg+mEebQmh2wOsLETWuZvsS9css9rIfxVheV3VHRgwdjCnceASO
WkZmTNRxLwA7T9hwjFzwKCNoKxXhjXEtnmWC3DXZYxbSQXfGdUmSpSau7k7mFX+iQSMpDlPx8XhM
LgDAX63W2DlOOsjIjHncuaIDy0Qjmr8JeLo336U8AZD0bDT/xFKm9a1PN70BNCIawnBlEqr/i/lb
gQMzxAbYPqL4Uzl2o8TSdRTwKg++MZt3wddfwuIOAxxAQkG+2hiL20Nq33CvtduZzaoRbctb/gyq
ZLU0n0JbhrrcR76xZFZ3KxcFCY1/IDeDbm6EukaxqiIN4hG+Aq31dVLDnQ2Dz8TVqNTUyEXjFBaK
66N9UzLyR2LjmRzxZFJnhXxaYoycUlvDLq/AQqr035+LqANFCpnlh8ZV6KCsE9/M5SX3rRenJMCZ
KiePdCPOCSZQUQzPCMGajptUZ0VCHiPuOupWFT57HH3vL+GOBz5YmKiV0N0dGYsGFXNvkBKq3KxO
t8sbhFnG2f+pXrPwhiI0LfYyeJU91Kjz+TlKqOcG149MLfgDB7+wi4siophm3EWerzM6ZJ5gfqV7
CRIRRWIQ8URVU2HdeWULZqCErGBzp2JlMDz26oRS+WVRf3K77pOmnPbvKzv3HHffIWvZhvH41iQt
J4UcWHsRyCHCrWYC+/1Pduwdt+Pf7HepOrs663jCGzfzr87nOjyEPPo50b9O/+WMAD27c7xkImng
aoOkjyDjn29JERCHNxk15FYsezptxi7c8uPQnHV+xKksz6SNMoiSEjS+Kv2KilmEr7zVsVpIoki8
Upx9fmLujobiw71hYgNov/Ok/nkE9wZ7JepwMHTFWlliAOR3BBuhB2GDzhKvkOi0cTw8jR/z1cs7
PukQpOyNZWVG0QnL4+bR699+qr/lKt5CMtC5ijcRU0SY2LFwzDH39PBWqi28oWjYArb5HK/1Q0aK
Z4v3TK0kVmYJ7TAE4Ikx9gnYFJvRjm/7iNojEPKJF9Eo2cdADsnUMRlcA0cXyA+J22aK40M5oXPz
+b+vTulhduBYG2wuDoCp/pxxH5Axx2JWAAyWtD8x+0kGRutezQENXZWoPRYbqCQ0vMg77f1+4gAj
g2/U5gRgYvxEJLlUl5YNRS/SpE8rWvpxC0694O4eeYS7EtwyyI4APo3NrOnxWF0E3xQO9SOnGUZ4
ePVfu4w/XMzpqAYV/2UcZOEaHE9rZNMRMLX9w9A/ZzHKGCF//Ue1gEhfB44fPoOaU9ssefDQV66x
seeeq4aJzjvkPrDJdK2klx2x3/0C0/jDQQiwgDDO41dQPkHohGBkyR0bIqhijwEWbTN42xm3MHOQ
0pLvt4dlvRsoXojQpDTjR5CbHLBfm7oY4sdEi1zBR5PYUW4UNthzwq6upHe9+kOzQdUPhQklKhX3
9Yx72WWtDLe5mgG9SnodN+lDW1I91/sNFswsE9AxnwNr9TndXbgPao++Yl9ZK/MhlIE1UVdgCMjj
VlZKRyaujc8jFQHPWOn6as5+9vklrn8ohZtw1iu1kE9rS7PJnA4R8K1NF8VOaJ3vOScX+2i06sOC
W9sypXmCTcciSV+lcdxqrUaP1NOh3GREbka6lad/9jjW2HO3xzwOX2vL9LtaaSBKsyG8czqlREJd
iuviaT5l00FSBswwaUf9B2z7jcqIXA2nTGO16hk0GxKNsn0TdAEbrkAq9dcxyxBWN5B+ivhpXF0t
/ltaxPMMZ3g80It7l2tlHtjGjMJ2BG2ryhFVC05O8gi/8+NMcnzTspYQva0qQjBm0dPzhKEGNFkI
dkH3P99S+2E/9cxnZQMEx2ZJb9OD8cyQrDWuGvxU8oB0u3rJKmU6Zg/Ih4a6zMwJXW0XxvN5/ydj
K3GCzVSxzRQ8rWgoOQ6I/iDw22tqzBPaPEP7mggZzxHxAaVolNM+Ylv1Li4G0HH1QzKH9q5UkYuG
NtdIsHGRtq3ykmn+opOYak26Q5fCwP2ue+wND4kA2Byswj35pzC+5vcEskE9KdvVJMAeGGYTVj9e
UsdkJ2rEnGLpONhI+bw9k9zNSvMOoUpDjCHitVad1MIWAb//05wUEX85h0tASZx5MA8NoLSNAwnv
t4ROp7Sn7X88FOvZ/twsmA5ohz9ftOe88xYFYf/Ip1IBP2JfStxqqCKaB7XBh/k2iMxkdMBwBDPO
7fkJbZ6pQ08fCFu48vef0ofJXN4CUyAyV3L52i8Pkv+i+D+L3PnHSriRGrUoJwf25JNMz7Jo4JNQ
0l0xZCkjvja2na9YdIxwdu/t1QMuR+M50y88N6Ifq7y1T1lmx0uIfH41SrxwdE6qTE/paK64W9pY
bNfe+1jdTJTj5wF2vaF5x5rXDbAYKD7v8RTIGJnL3v7Ir1TbCcUycLdjG1f7OwMmYD0phoO/rqR1
GSoO9NwHOtlhXldV7CZvRhIXO6HrzpUedq1fvEpX3NpRoL9BThGwNv2WZOF53EK8pr5NU8+0eCVX
D5dBePz1WztimCsyKN8k7L7/xqkaDwTBAAxvr8ZXrILXft4y6beAKttJRV4U6IjZmqJzblz9UclN
LN+4/hXngUUFU52j/IaF1ZJUpmDL/TWbKICKasuR7gb5E1IJFMzDFXhdmg1ilbb0aRONT9jHUhK2
ahbgqXrQkXWntg7cCoEwok+vcfk/KuzsbIb5GKld4+0w4b+35mVBVQLz3HNp6L1/CyJ5PP/0JvLO
hl1BbJPl9SQaGiN9MZ8lA3IQB5oEwVhBKWJRh3TjOKrHyQs79H5upJAlNhZau3MbFM+EuvVykNY7
k0LsrYdVte1jdBJg4QkyUUCa+vmya/+SjfWxxXKkAKvad6t7IJAYGc/7ny4txuldQx5aOaG1BI2d
+gecTM735Fb5Q+V3aAZppq5naVCUQz+CR4Tyr3yCF4lZJnf8x0w8RLrbK4CoSclLJI91FlDuo7rp
XTp6nKmC9t8/BC8nuNTdiMmN14XnHnpmaxdiU34KSJ6lRZ6YZJyo2sKOcWqr+A0Hl1KAykm2jq9A
pC67hY2Z1L2oOYREL21VfhgJnn8jfhinD+/Q6vsze/Bqy50unTRvuw4ExIGDXyPqCZHz/hJxO81T
ItSKPb0fQAo/rZLD2AWk2lAirAwm8B9fH3tWe9Hgf8mfxl+TvRA4k+pmh9guD+JTdNdXLC6xK8nX
M/LqD7/sFEXiPl0v2uD0+3Vjmv4PF4vECQegb3MS7ZC0alqXUB6xKjOQ+PvKN3DIrVN0m7pIUaQI
VrUwGY0EgkfqoE2dLC92tJ+vQzZpKxGALqeZEbIV6lzAUo0YrlPGbUEH7w03CEwFTRzGMdypblPs
YxUxW4fXUrr26fJptj47CSjz5MSEYgFQAr+KB18HRU5xTYeYeTDIb2u5XM29pllmD58dDi+GjiWZ
AucwCpX0IpN16tuL5IZOwizQ/xUbKXF+7xkxMYJD1IJcZMrHwBnZxJuM7pGIV2npcYMQJ6iWjtI5
hqKmgLIJRZ91QpKByxYV6lfWy/oCimqgA4kL+edNkOFfsowKgwW14hc1r2/gfbwohQPkx55ZpzJ8
Tro/ktWfk3mO3LqwFg0qP1PUxiN/5tE9GubTKWPCSu8J0YIgI910FyMgUtZOtlcTJCPhoMQs5HiV
U5NaLJJNwsBk8tsyY5HA4991HDaFAVTKHFnG6LdQ3DtLGb/ek1B72kVkHXQ7Ntm4Rp+2LFYo8k/v
5SmnpHavyMesrCZisBNf4PnpJY+Wf65sNxZj/Z93f8yWlwdvT01e3VSEJQp2fBzne0B1VvbAiCb3
UC0ry5IoNtcrxYo8ARzVVRnIvrvwqbY/O3NsVk82piIAGPB7qfQxU3a9DBtKkNYuNxan5ipel+5n
3OuuWeLPbwhk23xskM2Od1Q82HKPbAhpeL0aF4mXjJlnD+jILS3GS53v5jwAthmCWHqZyNH9G8YR
jjKTEBUFvb6nzBLfmHmSfj/HAef4jNHQXnv9YOl2pnmJuMVYsMfHhJIZ68EZCHmFWBnvIZHXDFLs
DjDqPNCK9NBJdMvQhXGnZY97VIj09HOWCU+uH7zUQpNdE96PJTYIKEGntpqLD37Wpi0M6paSCNWY
wLZFselR6VfPbBkqAXdPYxWnuRlCI9EcrP1xHi57DIxgFlDPl9rW+JSIueHnkrOssRV6UZm9CyJ/
VG7xeYCvmyjm8G9URkOyvwUnobBbu4Qghp+08r4ehPBP38q8nviPqxXa3qnG8a27FaG/rHvuurhT
rUIqdP3//t7pOwOO9vPfbMj7sJndGiBfazlY8t0W6qjefks4YjC6WqN406IOBlvCO49H34Wapjnj
VNDQsljwT23zqgpOzOIWCP4E76WvG/rUke1MpOSn7qE1mVlBLh86OO4Hc/POQ4WHAN61rHYUNWN1
hDQIN3kI9gqx9UcH1EAvW63ccH7uGtMGR36kO5U8qn3IMnQIYLMNnFRamqwtORGrJ5iA/7VgQWP3
mACCdRAbP00GAsQTfRh7jTtI0uRJLpkZk9nR+ArqwNcq+ZIIJg9PtiLo3SjTBNrTxzD7Xv4APC/f
DmocitSGA1nz8MYmj9cVv2OU3SQTh6x/Pl47iAoB6b1rMyAIBSVHScGlP1HrjzPkGnoESFN+qxGZ
TzNQjTXWne/7vv7Li1p60yuQLxqSwgQSItXAPMVQiyuJ6bFyI0AHdi8Zks/hFQK2i8BfCtOfCtHB
rf23K7JZ63HyrQ7Dw8I0+87wGqx8x/wCPRraeb9JZ+kdvwfiY2NbsmJHxpXBAzy99K3BtRwhIpA8
y4pwIhj5YXjc8Ud8piKen/3RukPt9Ur5xuKGMBggc45aF+KnUkuQzl94EUr7/xgUx++Jaa850hHJ
TIo+4fNhxjTr7UWF0alHYU0xDlwiBsXlwG1ggZAud+1PmyLmUwCgzXQhf46lJoDonW9xWj4xX7Bu
AmXYGOuKhqexMHhDgevi2Gj0Y+aZ7YoT18sxmJMFVboN9fykF59o1oLlAYxoIQJqBVu9RHYjuCmZ
h7GP/iEX4OG5By5oNE4SGYYgJCaI0W+6C/wkOFRRMmnMRWQG9dwXZycT1OFLSe62N2fSPSs0aXj7
jefVAa7Sl5GZ5IVfmd0NvOGBL3qpl2vqdrn2IpUPT4/+fM+FzBOk61dwgLaY+zVGxO5VmeTQ78GE
hzrdCyfOBQWS8IdV2HnPaXipDo8kVYgyxoPU00+Ph+IaL843vZTGlwzkzRvz8SDAI/nOKudhkISN
HGxwkJ4c3DN3/EcWPNKWXAgmqZMhynyyreD/53shBUAajpKWRVrFt16fWRhbFD98Cc07qdrLdGwV
oPiKdlIMkoQBe362dta/de48dD0mkLxIwVn3chUe3EuHzzdmcZpnEyTla1/W1iKlh9HxJc/ewVr8
8+Y5Sv5Y45x85bjxNjvTKN7CsWjMU/wfgggVcjAIeqG68SXsojQNOiI3QMG1T5Ty7xmSRdrkhD8N
ixoTJDhzZZtMgNXttvX+YIDApx3Rt8xN3mny8mjI95Vj6DIJDbrzZyXUfOIRJKupa6COoQvZTUPe
NsfzWquRBe3mVCd7+S/dtw/bHyysUgcw5k+rniqLI1vQk1dbg4nQrd5RSTPHmUbrk/ORSezmRxyA
djXwJeyDQHYpH6aMSTJcqjdi5j6BzdXTHnHBi8YH4z+Jvq6oypuyJuJTzDOygtIpJruSSHFJADix
afVXOOAIdCt0I+xzryokTdwNuzmWfKtrAlpz9fPJ/DM+dNFZILXLOmSDoGhTWh0Fhy4QZ+FD0KBy
in61aPavd1ZNTiSrsIcSDHZ2mvIkD0E3++07tW8taINzr8Zwdse9NhFKZcAi5USlylaTyBSPnm85
bnMRcshhdubJ7hBjkYsTc13RqDOA7Bd2aOR0QJrbZIBtSM2zEh2m/bCNztDso62uxSjB4JhacqqE
BxCCQxiiCFhtnJEkdjT/AvusWBQCGOeMGKmYVwGzqHZ4X1L5CZ2k5EsNJXpV2ibizZRay+hTT1pz
9R2RaK0u3LwGokHi/5xDHDKUqwy8onyr+933xPtaid2zmqF44PdGC8vl7IJAYKNfZbWtvUkZuFvD
vBp+kMc5nQdSD1WfzwB/9/IopIjwZUSEY/AjFZP7FuUdRjNNzbYjKvGk838ceNSf8V+aEt9rYrkw
NabyxHw0Jk/gSlpReenYva5lAPO2T0+NQXzQ1E8mEwE9XdveEuRvmOEFRlvih4SLvLKvMU8AVY4w
FThsVuYh7rZx8/rsXsTNLJIC5NoWZ3hOHrK/Wicy2aom4MXxQyRTG/lCtaaHpKmHuUDmrw/JRNKY
0xxNIOpP7n6SwWG6YsrLXlyAeHplRbe1pXD+BakDk8yeNb7X+sQkvDqvjd/1DSossNqsTbbovjNJ
9F4s7aq2Ldcvwn0VFj6OSsHDSdbWRf0DOo6dKW1sB6xTAWSZ4XKAgkUVm6xnPZU2VhyhPYMik4mx
FMON/jit2hJms3LNyDt7rp2mkAqobSscY4tNNRCCl1UqEGw6Ugqfn6Foq7HY3k/jetricuE6DsVh
DDHE4O99Mq3zL6dfSb57YpeYaEXwqBSzIMjFE2Yq5nMYLDcIqI34/4wwjeHbwmTYjtnNnJ/74UlK
hO8Z0P859/raz7yHL12MAWn0ijEjWMe7UPwJt0CKjLFvYscP4FrWW7E+U8opHMa4Vf9kKMVGtuQ9
8Z/KFivDjUkm/t+qJBxm0jUYz03ro4ClogCpVK4+iZSLVX6C0nIiRWnVEJycMlhpM1n9uDPq9ew/
5hU2ssr5JPF2Atf8wmlxmJrt4jf1eiKwkG8z37rtNlP0msrNcE4ix+fLkhKbV1NVeBFC5G1HIX83
frOS/X0KKvzG3NIoTSmooPlS/d4LBWnFc06i+FQBu/zgrM6fQVeV2eu0PijJCcNtOX8O0bpQ6NFG
dy94zd7o+cUpZmUzllGR3a5wz/YYDG5fAjl47hcKPIpyn61O6VXU1wVQi4XCnn0SNFr9+jN9P2kL
hFOZ3TQsh8FzE2uNq/fr5exNUV8YSXYGdRMNxkK6H2JDJDdk6fdvSb0wrYlQj+KLXbxOm5d58Bxr
jxRriVk6N2hxgtwTxDVt4e/PEmS23yQtx0oUuN5t3f/qdGdnRD+usKU4l9AnrtzoTSN/EQujTmre
GfRcdnmWy53DOOZz0QhTCpj8JJ14XqWTOLmMouC4OT9yBlTNaeN7S5CVy17f5K1Kx6CIx8PA0dsG
ANoyb0WKzFhez9qMpLLOwDXk7F+uIovVvo/3qyekIKa2RJpgxTLDleJGgZGBbstMxzORjNT7Lftg
wOVC4DRTwm1bBVqXBBcA0+tx68+i3FpVyTGaAfF+q+ahsmcJhb0VD0xq5pc3Y0KHIsjvg1gYpYxa
uzN2EL7TSxyGVq2kpvVlou+FvAMY9sLCwWWCRKdCbAKIfLiXdHjb6AV5dtM+NcPu4ZqYM95e5pVq
D4JcwflbXeSwmpFI9Pvtdd6iWhtyDE4XwroyhlmAUtWMSJKGNNV/GUdcmTUyMLSD0Zv1IA61UBQB
KlktA+fgX80tHnrfJchSdShXiudT4ZiJSbhRtX/bf0ohFpPXxHcdv+PtPslKqWGLwFZf4kyxNv3t
eX5IdoVja2abhljmEK/Vf2vVFJrRlbGeHhy3PRCNH5sI+mM/s8yAzoiAcwjTZhNMXramzdzJCqCh
q+p7Gxle/Pm7ZSd84b9KVRBqXSJunpAvPThphCFfUap8dr7MrxUIEkdjxvfGd0WP4KuC/reZvRbZ
XTMLE/52lDbHuj3bd1hCygh1Dm75r3PWQ71bFAEF+Par7nFPbooQmowmv+EKOeq5tMql+szEPJqt
n+yAYbFkDlp81SVzLj3o6/WeikWekCfxPDPqSvurKCXAsgoss9VPkaeBbf75etZaehZP6sf89s5J
nBh5uT65PhtKtYpPPFfzgjhE8rJjPU+BVaSpoEc8EtrPrU3yO6Adxs5Btwdy+w8Fu8AVqEOVnebX
2M8XPbRTWt/9p8XJD77zdVdS6mN6mj4cZGrei15Q/e61YEhiNqrLM4hFWAS1w7w8xMrUA2ZDsbv7
Kq44QQDe9mgf5E6PsASVFV+8k4V/1L8VBeNSw6NIQJSSx3mtNZcrqCi4gVAyxeoPQAwa/EICceU+
jXccDT80Gax92cglb5j682yiBTrVrAS9S3lYqmzE8MJQ3Bm6qXqndqkwjnU7ykxj5YPTcSjJzyU6
Ic+KA8SJ+ixt07CTgkUxvuEEtvj8e/e+Cy1xfkEnYbdFM5f+jNceEGmo3jJCf6hPxkOA8SHMKoBA
G2YLbvy7TpzXuJNAaSHoQzknxvNc1aoc2qF/3O6CqjUkAExifSTmFXaMFsLPQ9hwpo+9H2SJLoQ5
UGDs8+/Zj7vzWBC13eUq7G507SVaoCq7sCQxEWX/MqvzJ9TnpkiKea/IkEQS/bA0U5yFEabRB0xx
TFoCvyrePErjnfpbt5O1MWz5sat959SK1PyoEZ4XmwfT7tVjxXu6LFf40HfviHtNioKwmPJfTMOG
kgBr099Ue0wNFe9aRvRsC6OwDuT8jpEAGCCDU9Y75HoyMtTKwnTML+lMP1syRT2Jv+PdQF0dXvxh
ovrGkUxWNc1Lydr527SI3J4o/cXvDcDFXSCRyv9xJu1fAxC8yHdThlFUjetqlfN3TqD3FpBM+U3O
Awo3pbFr8FPWQE2UuNH9f8+MEV8b1Oup7zve1j02Lhxx7fLRWjpwSUkEdGMcJwEnPd00fqRb0DsF
/lpD/Shl70fPA/nUOXW7i5rIR98xDHbATfkkpx5i9IwWVbayjsnZ913oaH5f81BNrYOd8NbS5HVS
MtQjEus3On5+8bC6pxLS52pqBs0MaWMoqKKpVSA4ZsKjf2Ocef6co2Y7AlxoZiXUVGCs904kLzzG
jZgoY99j/v/Kt/OKflcbfJsjxSG4TAGL216AtaXFIW5EgUS1WYpiaxl7/pXztNRZNqdwyWSq+f71
Bwe5V+CDC0y8rX7K0NMaqCjitRPgb2Y+LGQ3so7ajhqe9R0oN6B3bPW2haWXaIfNH/2X5o6DkXrT
DzuX62l66Xqz+GDwE47qdZJ1ODOCsmldHMV1fc1lvJMhER2ApXJSG2AmafK8zgsl0fzuaDUoPCZs
JnDjQkufVkD8Pxw3iJCSRK8la7CpMMhme7+OR2DveoOH8RDdEXsxjlTRXrHGXbD2bfhlQQ9hFxSl
d6UJUA3dmPDvf2jE77lGkqIHM645QNkIJSBK0spgRn1/OdNVKjOf9ufnJwdy+4GaBrpnA4hTqal+
VBMl052y6knqrBumO+RkPqox9qxnlZQ6KUt4zltth/wXP/qdFuiJ2+NWyDCDIXQZWUn60Qw2Jtw3
cCPN7RzjlK3HmRxlgF8TKF/QbuPzbCCOfJYhxtekHg424v5lal86d9uH2WEyOE7kn2+VTShAYpiZ
N+OOeEp2xojhYhtlqBDvpwuS4Tce1Jsr7NtDdqTDKpyri0ZZ4yM2gyxqrBgrxAhIAoQESvE4xnQP
iNnn/HkJ3ufrHfdj4/YWrMimEIS7nMbFFeSNVb8J2ezuftxIS/zBss3/d3EJsMJwN3LQBLJdjiBt
MbuKTbI/zzQPTV7O48y/UcrJ/GakG30zdP5VR2yGPVlTjPbN8WfN0DHCki3MA5SnpRKIr4RkIckF
6QPadAJNRfUkbRv4jMupfxzJeOu24FIiwczOGN76WkntJRU5BbFQKgVkC+l/CBC7qbLPNPZJZDYP
mwL26QbpLbUBEfm4mgknb9tw6dEVstcCUmTqzuUs4TXx3flUQM60om1XpRB4NeJEegLGErh90gkh
ZVVn8mtmrqRaZvtY1zsDozjypx4FvG4jSAVMjnpbYEOS0otZoA4U/jVUaW1uxspSlX5Qdkgv5KB6
N+/MOogtPtCpgxGxCKocaYqGzZ+bidCOgNCLsTr1O4qHd3SURwZZckRAQcU8cpkfmou51PeKHO42
C2YutP9fmis9cEE628mHtKCppsI1hmb9pNgU36wx8BBl5xhiprl6lwRl974ceWe/to8eVIBt7hlq
dyYuXWRRe1RWqtPXACYnFkMHo6tTj2Nvf9cfJy+43ZOoVbMJXK2oFgy/W0mk0apA27QXEm/k9Dxa
/kCt3LmNshOZT4iJDVs8VyqU1NJkUn3bLk3M8mPjydVPfBYeZ6IebHn5KdfTE/cceoCFjv6qDz7P
H4/S7pFVPEOapv9camDrjvi/bJX31XtorWYdF2R0YasP3y0gxqX7cnFD5vV8srgBTkdb1e4flS9p
bvzDcrYJWV1fCaWILKJiniETMlLpJ8Ps6LhgVskNhrWHp/BS6vGrpx5D6rbfKNpn40ajYTvmGnws
tOONoV1Qsponoi2xZyg1DWjrs75AuEmFMKshXoGnGSE7Ukxv8ZZzUIhC6ROzAZarY8xEVZMSkyi7
zE38r/LDazW8I/R6dAXblipPDk1MbSod59Bn5q1ec/0OfPNRpM9S7t7FqnTpqwlxl3KXd9FeZ8rw
JgS6Dx3qPRRHAEHiWNysmAgrHWb7VTd2otkaRGz5SBSfqyE/swIcdP01f0ZfFMDXiXzEKgHbeJwO
tvTyQMYlAWpqAvbYRhVtEC4DMBIzkhxeGqqpNFXaKA9dERY3Pkd4dOclse7eOZ6U0YWaPj/IAhdd
jExyqVaV8NhRfli1zOwfjYXSD2lEWBe/qFlyf+rqnn9eYEzfgPYrannRIz+eB734RwtzsLrH1h7P
g3s3ggzOEGqXiwgkxMrvN/3nmDsohZ40aozzOr6UmFUPZsSzmAlbDidIo5OLeQeE4DzH9YongxVz
cf8o1l0jmNcf9Li3qBDjfOOg+HS5ro+8yO3tk5f2xRLrmeYTCcpxsh/JqdpTrpLulPYEbzLmEvay
iEVRZi6pJoqBSIE5Sd5d+PWZLjXZbRFjF00H4ZgDPBZ6MStJlM0yz+q39dgA5ErJGCaNl3OgbekS
6yFJGajLfK9lJQcpcKxd9/rO0VQ82YkfBIWd1KGOZssT2gBLkN7KrFtVCvqZuW8klNycnDybu5V/
D67O6fFkbiA/YCGqqs2I8z/r8Ec/Uuk5ANoJFVv75ORvFXZO2BhEWHqeAsli78cjaKgzOpaQKC/V
5nfV4dKi5gL/Dg8lrr4GuKDVzJu91iSJEwaxTSorLm6VMPKI5Izu7sOS62Fzngc/hOZ0dAYpNmxI
SEE9ONy/YzkrNHPhb9OokWeYagcXzEys0JSGw045THm8NFtPIOwU2qb0/whqp0LNIQvCmoIOUjY4
cOzAvktKZe5Q9M65sCB1wD1FglcMLMKVwEoiDIM5EMiGq0o7dCTnwfbyJiJqH582db2LV/GpNz20
0H6tDF9r6cMQFkAif80rF+GIUxTHXv32SyxmykUdpBmeQaGjLpyFeMGTbrDrSy2IYMipo0s9Nju4
G5rCwg1gXrKfCyR1ASRBK2GD0eWZfBy2aL0gE+G3pxtqLFyDejV1FLRod0203zQQT9rXvk7hWyE3
YnMf8uRwCl3+PyNqnW1XTutnQyskRxctZ7PHfJaPbOpifZgem3uACnMPY4rBxp8Xj8VUeivpkBFZ
Qm/ajMHEeTu4ggmYCN6r6A47b9S7DnClArRvBdT66ASj+PTvHC033lMbKAxL5R8xjpUKA0ea6NaK
wcMI74QzNV8ePIW3BPpdhmdweWRJkRDQc/g15v+8ctcHfEcf6Gv1f7OdYU88iI+Qh1TTsm+c4Aep
MIAp/pNtRffiJ6EXzTt14btjVQ5VAsxhOCFuu96HlDL75Ia5t7syT3YctsFrfiPiqxi7f+ZGpwii
PFg5z/LHpsUQCNfRNoc1Qfo+PvWcQ0S08K6J1AYttbBoUQd2gvEmQYtLqPa/rUWBeNcVcWZbq28C
mEjoBWLaM6AZno2zfwZLvrCwiLITMdqRAPSJX1FADourR5umqbZdCWX5NqDrJBHRL7dgy0CKFHBc
Dpkp7GTPsyJJyjlj+rBYVMPydPVtdU8u7/z4/QJ19fgx9PJFsj9XDxWXaFH9oPHOOKGrFfnRU8FS
IztIyrUjegW1JFZbN6gOiqKIYgll5tMqT30e7by4E80SEX4cQ5T6I4soc5NneQWnLMtDAZXWVfWv
ml7MA6aFjMoIuds9dn8sLym1BHyN+j4VsX4pyXgWjN7nkdBeqEnndICuMrdVy4plj/8Q6m522553
CxjnuuJMXdNRP6fge1gA2xEQ4x2bD6+YMVY2XpBgQQXi3zMs/7OuM5USUuReLleYRlLnBbhpxM6a
Y/8FR3PkrxRkl/Hi45bD92oTudOGgfC4Un8I97FdY02WMz4446YpsoTpc4v4NhBqr9Nkpkpd1df9
Lh2bnwQMSCQ3qZTgHQojav3wK5wPwTJ7b25DXAtxoVNzjZffqjg3P07EUjUnOgUjqrvFhlnRtRKO
zjQeU3tjlkg1XnTRfv0+PQjaIaD18mggWzr0WH8VQQ6aJRW/jdsOEQ2wL0BnqYfXLqF0DreyJ30J
oMbdbwvQQI0PKPXbx5CYNYDm4lsiIhjf03rQQyYCI5Nj3Uoxh9b+otMKl/FkVFfd8YRlj47i2hJA
0LsHToWvrfjfyLam/mWLIAcP35WHDSHvLuJpYTbQa929hMiNhyBZMfiTOSNtBF2J+XRwph87KbAv
f9MRcK1PtvL/H70nrIs+pcn6knbHgw77GGSMdrNQgW6iUTTIDGl+ZYDhZ9vLtzszyS07DfkOK1RU
eL7EIVAUwQK5jRmdcp7fijEMk8xBCfs+mbgSPJ6OHQMpmnyYhy8Y3gesj3irh0Yn8+A/KxSIGLTI
SiECp+Wpm/iK5bdcoojzE/BuJl0e2E27xRHB+lAid4Y8FhTr0+2dAPwGhjGtQNyhgLFwKVkWWCia
bt/mSettTw3P82vIx+PI5XHRTWo+S1B7SslRyoG7vwBHJd0Y8URHVlnJ7FfVFR9ORxFvpTg/bnH4
24uNjdLUz5sK9Hf2y+nIU32RhX7dTjsnKJMC7ELbNRYMJaO9stSqk7MOt5hsEwkuFzD6QDVp0fqc
E4ihRCCrvGjIs5bFMJWtINAJpEEYo6D9qkW6IwHnJDwE4QouF787a5AzHCu6Dm8hz9bs7QNnLvOb
K3TTo3gdDvTzrKw7w1Vnh3PXXX/9sxneKGMyYGSK53x/MIw1MB3K3T21bNeUdni+zoESLy5E9PbJ
Aoh9nfTH5qT20HFe2OcLHSMsEDGM377gx329I28eJEFgz7LNC1OXbP2vMePSilqj/QAmJecdOBBF
UXpyBXDFcwq8P5UauPn4UHfBh34lMiohU/KjdkZl9YBwpTeEHP9dzaEGeezDGbdUo+Sn/+mSIjXo
XQFWv1+nteWpkWAHs1/I5YsCWb/kefMSaBWPPiAcWLnzesouMdrL/Blu1p1w2hMyD9X7b2XeP9J7
Po5X4DQ/GQ3MTdVDirxgq0RT0jWmLGYSOq3QQ+SPQrryE5tqjMxEVeuPiE0snH+2hCUKSQN2nKF4
S/qaxqbuEDopKTkiNDx5aH0XrL/G9usgctUixOR9pb2jiVvrFbuCtQBFXrqC5i5KN590E6sStnz8
sGfdNOBzl6r/UcNy5g9kCPjCrXEaadmmyaY6F8WzvvyCBleW8wJRqrEA+pZ95p2ReP2fjP7gal00
lA/SgF1J6BxWgPxqUwKIhpIPf6XuA9tnmm7G+XQOvL+7lPS5neDFcimzQR9KOlObs/rUJFJ7q/Yy
GP2K1ZnUkOgndUlOLH93oE67RvLeHXjM9z7lSSTxP1At6PakFigRyzVBpGfNwt/Vs2ty6xJeTMXh
Uy/466hybIju23GDBi51hBZ2wvJbhiaDs1ah+noUXy5VUc/oWJlEwaOcccMXzgHQZtQY+2uIZKNN
bG3jUgCZmBc467ljB4tJnHu16YXjHm68Mtvz2IwS1zgqItsa9Bk+A8MurA/0WaOtjHNaI2U3xuDr
ENVnDnDwhYXpjFXMNEE8t2JTKcoWxgR4cNVcsACfExEFSYA07jp0nqEW5pUkK9aCRxQkW0JH7Tea
ZHrm3r84X0ooN8wgTpXqHtHMzdnZC2aLS2WVgpzl0PNiczjjW3+Nf9Mv+QRjqCAWjPRrNMqPlRnp
D/vAJePHHDqpRRrtTYKN6qkUq7srb4ucAbYPpc+/4E6V5nQTc+zulk6Y3bkgkbgMYZ8o/ki8RWo5
NvSDEDFhjgi2MuZmYQmQbT3ExWdIE2yCk51D8tRtUJvoash/2HxItZwgdgRJ+/nDc7TnBxMmfkck
sAPSJK8bbmR6Qa1gYIClxtdJjTPM1nfTenCTIP2gJiL45xkLIQ00nI9bzp2YCs773iu/vbBf+ge1
EJu2L9W9nC7zqtvPPU+/8/dQUDhLRTgg9EiTAQeCUYSopq61gKgA8Gm8eRAgqVIdCNLEmcZMCk3z
0tRvXIbmiqy8wUQXi3mWZJgpRm0pBSvZWBziaNGRaT+qRNfS2OQr70ykIcT9qwdcsVcMAScmAbRu
MxDFT9g1JQOhO0WacdaDk/41YAAxTtfKUo3q9GalxYeyqPc6hf1E8xZkVo11eNCusDYFxBMKrnCa
AW13QkIcidCZLAEIZpH1ozY7DRIld8trc0Wk+gntpsoM7BdGdrFf7+MB+f1dfy4VTUCXzLfjZFH5
LarCBZlMQ4+tDcB9MVmCJD+aMMdL9Bxi7kS5YOf+R6QNJWluk6ICmkk8UIdklg==
`protect end_protected
