`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hRIovrUsnBxBXUuLxVRS+mJ6gjQTWU5BgnftL7AlUpCi+oDsfKiA2dBlt20d8vRSmxzZq6htzycX
O325Y2lVAA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kBl9IdCIM3o3Ki+q2JZ5+BFjr679Xv+VcTquxmCaeCn32y3hfdQdmARjalK3OvJ0Yp+fFlA+rOlf
ia6zlEba7A8ixmZBOhvgpFy+epsIMarvXQk/DgDU2mlWi0tgSbBMHckaG7XEzdnYgK7yUgniJXbW
95iGCd1eHumcPV7nL8Y=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rMTI4EPuGy+XRyQvnouX+OUf9hPjA9cf7RYlXSDOSVku5bMEPyC4N4o7Odl7kwNYb80HsMgDd4EF
Lt7Zb/Z6WOSipNVP9Gf0I8gCz6hf4jNk/hVItZlgCHueVWrCemidbHTvrYBaQdzccA4qVXPYIXg7
v5AGiPv4AeHkWeBRF6Q=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wYI8P91BXQv8F7FCMW12ea5EiOrkEtcQMiYRgeKY2xTCszunB2zyrlpwrZw/Jt91uMSdzgqyXFUc
FA7eZPY46UU3bQzTowpkuDMY9TwMGOmoKABaPnO1l7W/PRnFyNHIYnSfZU/Esx2qoROUGW0HzovV
jM10c7eRuA/sYt8hQJpc+4tTX2qZkcLNJllFuN9nOknZ3pJcUnjqJf1UR69ySyUNH2ljDIa9KkVm
JTVkFeSQPNrFruhWOqVXNHOLvBLJocnrkykem+R+SyGEw6uEFlVR1HFygSlk8djVaXZlxZ4CVBkz
bS4Cix+XFQoP3HuIMDiwRskpb8Dz0hYMzV8rXA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XJs/oLDTJq4I7uFnRGdtD71df20/IhUx6yiZMT2TdyEIiQDiGwpZwBz59npVbSgvBrEN9aSwt1CT
3Tga3nsAm+OIsfMy7cfW9Wk9T5be5cYWmRUo0vuc6+QVHFh/lr9K3F0A7wHZALhdPR1XNLSPzH23
EGCBLdyconZUaIvucxBbnsnYbZWUnu0NGr01ljwIbuOjZNjkIhtMR69xxaC1YH4Tfrehq8gnxLw7
wM2mpqeyOkty1QxUzhT2VCuG4dEak6PW6PWGx30/odA6Drw95vNErfzUrqlQtEeDdm6Bw1YNr8k1
8iIw3u3x6UO7i63Ke33Nsw10TRNwcjCsHlwl0w==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ER2HyVPWy0Q/7TG8rQ8YfAgM47hJSBvwR1ElX/OsHwyVFv9BvfQrcZLpVRxdvxmGjm454/KHu59l
RA7LLZBzuSLwPvjJXqEMMnfuqTOWE8CoeO8160Oe898UJIIUt7jycJQzjxHmyUv+8vVQEWE3xRSm
xutQbXkb+FdMQsR0+1R/rP8YqIyjGO+DqWGmx/4WKP3r/yBQW0+cGBDSx7Q3w55VEnbOA3WMglc6
4MksecD/85SwcJRrdR5ILZnjLq8GTZUOLax6BSZKAirUsjoZeflBscgwr0GqE1VSxmXQwnaKeP4j
FrV46LgwtuGpgi2qmc1sMfMrj+ZAwAkAMJkMcA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6768)
`protect data_block
sTFPVpGpXtoBd+cMsjynHfHug9c9VAJ4pNpFHv7gDyjnXLchUck/V7p/xv+QcwyAEQcU9fi9CeX/
IJND6RjZiKkcnZ2qAMf4UiuLSnPokcHNNuHtmTk/auiAmfFrIg9B7cBDf9tvV9FPxHpAeDcLUZec
r/KiWuWcK3+jnPMzlcyLX7p3dmKnY+MlMbHziqftnzkfhVMjwLp+AV7stb6LSZSTiaCN5RYqHUFS
mbXyfG9yiEDKvqck694lLSeWJaMtkxUrWkcz4eBP0LE+7/fB3g/CQM3J1+bzmm+GIV4WgH6M3s8y
OMpN7gVsTi+kpnlX6pwGwc7UNUku42KdAh74QKSeSTmkQH0GzapjMPBLX4J16aCLAlG69G5XL72u
X1PTxxdwcJypAMpFQj1zHgv5z/Y7Bkdbg5RIeeoBx+KzVsX8SnyM/vk/degRrBAsS4CyeYrP/1V0
8X1qtn7bCwG4ZESkUshQxqqYQzlIBnyFLWr1s7Ksyywbt2xNEWSegA++wgsnL718Yn4mBku3W8Bq
L2Gd/s/dDxEJlE0A5sWxkaOqA5t6nWCPSsiFVp+8qq/7sIeswUoTrDunM2dyTtw3zhhFDfaPMQQJ
VpHvZ2DEVMaFiMllfRcgru3KZ1h9wuOB+kFSs4wByRg6sFEQfun1xyWz+zwSNQhgalw2/MKzjfng
tx2B92tTx+LcNC/AlfGnHeYIWNqcr5OCPQEd7CoaUy0I3+/amqErLl4FgYmFhgeJfDNxaGlzd5+l
ReSR5Y9HnnWYZA9gYREwK8R12zmPW/Wshzh/wK+r3uhwINNL1+yTbInoZpNvXUj6QdMJcUAXID0q
OZRGNlAnNi/zWDHWuZ6wVx18nR8u+NTcNO2RIN0Jm0gLzcvaYxYokfaS3tBD08M6ImIiJdi9X9cL
A//7JyECbJE/NyIzhYILEWYVAcSyjWEb0X6upIObmzih2sWNn2Q0GOcs/e+9g/L97ZlAV2O+SoUY
vvkrrrP5nLQItn6cAWJHVddD015I3U7zylEw2DHgQ6NC5cS0gK4SapppbJawlFApmu7wIZ24Qw+z
xFMTqyAOwHxafQfSCo+VJIt2xDPYcN7B1eagPv43/tcL/eZbpve0wRKcGFxsXT4FcMHo/mKBRXft
6yfZU5uVxYT52VC/zPgG+E0PjJVauOcLcaFsY4YyqvEbohEJZ1SkUlWpU8kctpGvL4OoHLjVYJEM
NrM87P3PCTe9BkqGH0vv7POgi/VwGbryrio1Vt7KzQXbzbIThGmHWOcHK+XvVjBhqsrabqgOyb9R
38fp8vOZwsTV00WkcPdgoPx7yX8146SDJzscB4+mJxhTcF71R8Rk+Fd1UpizClaBMmlUEkoo0Wuj
hzPYrbLmWet7+twMw4TotXZA+RneazndlH+66jitv4mTHuIZ+5C8oOFXMFL9IgkicoxfzP8vm5XU
oOpz+EsN/Eq3ftV/TsnVQDIkT1W1ja9VnrcotmM8oH20XwAe4p1PM4H7Y3B4NbhfHglzrYfbp20K
3iErev4hf1tiF4tGnPzQ0f95JK7m2ppJmrXQ1y7ylgJbgq9bgsC0YttE3saXfTZ0ctkCg+IOc8RR
qRUIm9MsmmEgZZ6Mv5xWpV5BA8wy6WOl3i2XIGtMs32sm1biDI4U0JzGjRBrBKzOp88LjEEKvDi3
5Sb0MObc/V7CYuUnVOgxHUSMjF/YmLORKQJ8V/ca6LIXtfAh72SucvyoOyjw11t5VDgJHh+eD+AJ
LCp66CvFk3rGDUx+VBiWmExgNA3koDWaKbj0aK/iO3sx02AuxQZxon7lrVUKW2B0DYT6675lmqjo
ELkvxq5Tkthw9Xwdow1HkDhj2raeVnx9hWesG+u5NWYFW+5kc2xeq5O9aFCAKsZ89cBDJ5C/dhMb
k6zgc9sJ/9/gcw8gZjdHAbLpQQFhynL8Y+XzLxOaaWTQ62SiTzs0jQOq4dVLL8Rl8JhPDW7usoQg
4cTQ6/sKm105ke6ShTRZsodG6NTwwrLw8Jg2jcKDWnTcR+ivrH9zEDrs8qXFaAfZPKf0js3UXfH7
iJTUPRc0IdZFeeML+bfvpi76EDpgXefuu6mn2jk5l2XqVyXiV/+rAAtp/eh3T1ExEqNjTMN5Ptjq
LFLr79dOJKQhWoSA0lOBxStxrPKJOW8uFsw6HoY4z8sTBGSF/98sJAsBIXaRpABRQciOXslzYPNi
shGVjq3GATk/NnAN+q5UAWyAW60RtY15KQSZm1JJHmp3xY3zeudCDkK9tEB8nvDgjip22nX223p+
gVlnasgsplbKN8Y+p3zCGZEDkfHyxXnW3GAHB0zMRJohrTf2fITHx+a2Pg1duGYlMa7ngCy6yXYP
H3MHrZIjXpZWKwBysb+Ih9rc8vstH15A61frMJiVXFSikRxckP0GCvRKvY70HyFqs5NcnhqJu6pH
fdB5hasIX6qJF1Oc4k1vbRAjPsp6cyOVBzcOdkw0ABEBA6jdouZVUoJ8XOTf7GccMZD7I8Kb+44R
mIDlgRltnWZV8bZMH+buyYJ1K/x7mtaFEkwppJg1ou9VZNwmkMiZ6CP+Je+Qzb4h1xnFUesKveh5
T7jcrK23lIWlt64EFYrZOCoaxVmdmXyuIecPJecCsAVq8cz0Dp8461MEb7A1tjhKdBa+FuejdmLP
DkihzHka5jwOkPbZ2DchAlNdyktOWD7GcPmH4U8g/2cuzcRHEVK4VfhF9tEL2GFjFmGv5gzZFJOR
Ujya8RNLIiuVA/oI9P717pz7T8GLTjrQ6g38hqxyu58NoSxEMBZcFfuMkWKrTKSxv+WQvavLFJ5F
dD50H0EONgMAFkVdQrO9R1F+z5J/rJRWXB9yQHq4Bq2tgRnqk6zBd1zPKsA4nUXAXTmZAMj9i6Qc
mq3qKUfGS1XCV9Yn0WEA8MWEYYvwjsvs6K3uusHUPnnH/DLWV/EYcwl+yO8qXgNXvOsP5JB0bCx6
DedLjaj1+E+4uDKfdwM5q4h0jRL18Crcf4lK54gYHC1tb5UGA10WAzIsh9m/eenJmPcFIZCkieIc
bwbbQGy/1MdyCmH5FXlqztIe0VL6dx5qQCxW8Z8V3+u1eJyO2yLG2Qf1IPz8VhFqLIjNcMyTVqLf
AM4ssTh2SGxVMhJy4hOU7F5sQsDWeWlaoVICSg5spBwLEMkJ1pnt7amzScnz+kCVkEoovVOS/N0k
c8S4tq6he8JhN7x7QYBM7YKRK2foz8afFjXCu0rHRkB3IXrzEMs78hUZNN5KMxS3VCyqC2sVqPAq
JNGyIjmd0R1Uj1horGY8g1ZaAISTwabhYEl769Ltju526nP8pf1SvKDQ7xxAxQukb11apSPYVUHX
ik+rS8TZ/DoFUndNvGzM4VmQ7ixFf8gTOnpRnuv9K1g20i9DZDYABldHRS+MPxqQtBptNpiiF8RV
xjNtvBysPDNZdenO8my9ImcPiVo+p/qbvbDISrazYKOF1ldWsU+9Z6YO0A+qRqHlX5zL5GSLcG2b
5ErsbmbQVeW39PQfNpf0NYvvTLo4wcRbO0ZREnpvJCffFjyRlMa2EAeQ9GPs/8nExuYtmfr9U+v7
qBxrcad8b8FhC6Dh8A9zuSKFDD0GAeRdSOurjutiaq5lfSs1nUyjjEFbjYBpin3xMtm40Fl1WUwT
jXIwzrYG0j5jklF7nj5FnUeYdBw7eMP7H/CANIzK3X5n9HDjHcwupYkbC73PQgw4BVn0+pNPnUfL
yQUYp4RYv1CLe/vO3OFlP+5bZUe3EbGJKQjpHvhEuxZgWlYdnJ5lKZ2aQx1UX4w5Di6flr82Jgd+
//hVnIyHLPTtpOzx+bye+ZjH+zD8ZNPRnaSo4OqixGKkh+mf7C6XiArhaYLmcNUd0DEUcygoLVXC
gOYJDgb6rJb6Qp5OXSZEgUf2t/l0Wh8INr+xUZzU938auql00pu5HhGR2hKIOijcfQGIL3wRJFas
p15OG0T7qPGGaZyiF5QSCcqVS0AxmySkqiHqqGVcBDQDs+1cX0tZ03HCRWSPBa6bGeUSZGcxWxZY
CJFwrMLZGgjs9zsEMRVVijgC2p07hS1V2ySKMXNhJ1Z0rzrDO5XjXE6yN+fC4m3jy1/mRjy/vsU3
VdxRrLqMaEJ+JyWxdaOu8Wn2TERny6oNlyQE+AW0bPrX7JxNy74v9JEZiPgLb+A8XVcXCJsaPBKZ
eh/txkZkPupxPdhNLyTtwyRaWd1YjOoJEqvilFhq11YYcT87wW2n8w+DlQYk+e/423DfpvkRKDCz
teiFfJBoCstD7uYtPPFtWeUqP5jmZwD87IZbOf4bntiLeKMFN7TCYqNPjzPBwLzugT5JuaRBz7BP
YFfVvybDCHn5W7YOaV+way8HUkMY15+5aKqo6TEQqesuXhpWIcdAY/MeaehK//YOKRNrhstrFD4/
sw+gCKj0SJjYePBAMHBf5XvmaCSUiECxcSBQQyEBPOcosgS/iFfY5l4rqKQvWZ8TWeXzmYwSATXr
8azQD8kizZHzOmcwjIq41Q1znHGN4CxlQuxqy86PuGMHP71JZG3o04OGjDGjdivlCUez9HPxX9qq
Vvmf955EpGKIM37qdhDU09pBGbs/D5G2y3GTNRqq2jaNquRJoJ+T/nknTw4gz5/c23eOoXoxx0ZW
gHVthm5FtseA+64ZC9EdVYlM6zU7XVz63Z9ZYB+RP3+xXIw+ldadLoonHmEOucbUtj+XYLzFNfhC
RR8ev7zFfONNXXHPXGG1cY4OrC04K6BVFohl4k0D5xKkByt6rprQeUMpTsPhECvEJT+pgkgLE/w1
b8WvmITM/tVG41lPtxsppiUPqqpetSpfbSN+4qsy3QK8PUOFX4jmf61nqd6Y4whnHExKqAP8/43a
DcoJGs4UyK6BM6hR2bsDxjbi6A974Hc/4z8Y2iy2desn7Z4ACM74PqrDRFwtEifAA6Kptr+JlvgO
OV7oDsR3mI7VAtqSKeOr33sk6vLeCD2MOX1IiIP+0JrCTkBqetFJyw4v2jvhYezeYLaY2k7lIY5q
4d0CNG8fxG3sJ478cDAW5tSo5/ydmqgnsOwGlEacyp/0G9etd3Y2H8NvPfCF06IUR3954SGDPQ05
wNY85DVaF6fVWXZz/DrbeQTzmagmFnjopa0D2To5TUcvuMtzLwBzI/JGdx+QiRa1sNaHHgRqbrIu
ZYEgpO5drAHwzKpxdQNTRn3CUq+dxqQneDhE2bGSj4zaVvEBKePfOO1rmCsXSq+mG9lIFnCXQ3Qs
SclwGEngsrgXyIoXKLeR7pcpqYdwEThPj6hJF/Ba+rjjMvPQRxwQluao+YR23/pAv2ACEGU+VpK7
ZllTvUCTESRNn06lptnDEu708fj1HXC+a1l0R0+x2q38i+0bmHUztBBUdUgXMRs9GQVZBmJdaG7m
f49YuFQgMxCaIGkqzKqxvYW1bjra42BuJHH7rfmC9f4mEC1zGwTQIEF+Ds0Z3p94752pM+wY0g90
06+bK0pzA5XgFUBObeCkBmBX+jOMODMwPI28gHWhbg2dowg3yZj+960uDV7sDnYbeNo3pRAfPYvk
r27777vlocXsP63QhkOdrtEcQNNYRVOf3W5KJGnDcCLN2tAkoq/3ZHQCHkMbim+Du1ZkEn2KRWgc
vFIObUDCaZjNWyOzthVMdKFwil4q7+EAkv0mDqr5Mq2uSxhZYw7CAfCT0Ebtn4cw6BcVoyHBjwuz
CSNbKyHqw3F37vIUtcRragMGSfLkCP/Abi+BEAgVoFO36gzyEHhNnIUytYUGGLG6u5xLbEs6qJhr
+q4ZM7WKYq008ETz/uMbOoopSJMxCnXwc9XH0Z3XFarGVaicTQIGQaAoQhduU3PiSwGleyhz8zLC
X2lYPSKs9XCZ1/Sr1piFYBBg7Rul5x1o90iUHii4kM67EpTsliY5wZBYFbMPZgkE0uJ+6DH9BeVk
1mzGSecIxt7CRdXClSxBSSQUFXGp6AQqG4xV4ZwYQU0uYY7CTuIUAtZhFn8RG4R8S9UMHqg0tvQO
g7HAfVCAlHc8lT+PZP0iQ558DfqnjV2QiN9Jq9zT67WxEmrJUa6ypLcdJXO64yYQK5yEkdTNEMeH
EHLTmUBn5wNdrzTyZMI9kyyTakgPu8UJicOpiFLMYYiR0MFDPjFh2GF5i3wnvazCTn0HdkmXzdj/
cxk2TeIBrRCqcfe5Yia6qIniHIXUoEDt36bNo14AhC2JGYV6kJ0eeQ4bOBnj0mCpiDwMtm8PQrqS
qg1dZYONT41PZhydAwmd6ES5KwxID4/GKjLltMSYKe6qx8sFdKqA99j5cZA5C3cBGUMcU9sOrqpg
bOQ7KZwW0CQ9nq6kt5QeROTbv8rSBzjzQ4Th5KyY5tMTpm6n9o1LmOlqlJISDona0phNnDMsXXeK
k0hbIEJnDGtuv+iW1uvBxGQtjnJR3CBtyWtVw/yshx8LlZjtiAIJdAmi9nY2gg+DJOIs235hDXx3
sUtxKn+2L+lJe7bX0HzC85nbKo0HGuNcbCBnYtWKUTbYqVW758USpQZrHoXCps7s/BMftXS0XMHM
uSH4W0YRB0lkW9aQSldgutWTfDVxsr0t8ao8Z6Dpgf8nvMvwSKMgV4M62rZHU6q43EtBqKY/O+Al
RlzG7Sf+hm/UxfHfzViYlJK4ShVT0gSyyOZkDoDsUhWSfDQKQG65u5gZ1H807peZyz2Ph5KyuED3
G/1nBFxPEncrVslZ9bvAYP9zEnvijzsAhbT5V/PE2cwIZOooL8RGraLQ/HlQw3DdRT3r6bzbAlJS
J5dMdjZnRkahsfe+TP/acMrzrgHuMmXWqWx5y2CDRcflzsr+ei/7Cmet58YyohX92vCpGfUIaJON
6rz4PVLN/blo0BVHO6Rai8OVJrvFuBtWXsnYdpE7wK0cQuKshRchZZOgi+qRiOfdeCYuB6Jg8lQH
aat0ResAamN+Fa4Ka8uy1uXTD+3RNfeB0j9IAvhwJz2Xio5tjD9wt+35XDLZId/tWsi8oHKi1d/K
CeimNASnxJHpqRqqZcpExgOM9mph+OZhslBR+hpr++WlV7+j/diT3V1LRJ8/S1FsryMfEurMmkBl
exZeUr3AsGcXj8dXWsQF1SFHe+B+F/ycSYkIu2NgTD/gvaqfJRzTVouu6IgppVDA8yFwU84+fQAn
LYzZtqnPAHDbLXbhm3OeIP8EMFV8ws6QheVdQQ3aFH3Rhmqsfsjth+p7Q7DCZA/hZ3GLMfTLb27N
ayI9yhMDod2c9Mk4oS+iRJxXYOpnZT/ePiSA+ESmp2MjJKxWoQ8Gl5QuX8m9sCHcQtSJt9ifejug
OlPj93b/UYXn2NUtLTc8mxXjhV5o9xq+M+EAvdqWmTJ+yl33I2SJGmjIh19cz1OcfNSODhpGrleb
wRAGarMpsk4KE+ntS+EnYVXA/r/73gkvTHCXC+sYbc7beoIwnZvsvhDwxC+Jep8K81C3/yeiq2KZ
16fofV8JKySezSqU3mkvKnDWZ+Qhphl9Vurr+HcophSrKWofDCCDqTMC9SwH84/xZNHBWq7cLYqP
9K1dhv/QodQFhPiZFKTy/phcBXWPkbcWCD3YJjtyH+8i6nFdbjqM0d/G8VpL1LVuPKwgtEvQde19
O2o1bGbrEYOaQmvFYNnBhMPp1VMTCTu+m0Pi+XWMqflFjL/ediysOEsm6HanskTDDYn8qlg/MW3Q
pWJg3HuY8eHhjBxHE5hKl+eFu3GhNx4meHDSqbBybpxoczqSZUDfBF6lWoDfvHFUOo+fPWbz0UMB
81QuUGTTH9Mu/sZ/nPvu9kh5xFXasVctSjAD4MjF4x+Kiz0FvWS546a36nBiwU/krZZEb/tZI59h
gmtLnylWH72UzauRPBZQXj8HWPSSmQkkyYYKR+56wa1t9JP3YobTZGgL5XCS5jzgIe3QU/qZu2u7
6+gZ4ZvMYpDPJmumERoV35lyiAfT7GM8qMXEzBcdTzwo7V7rGTFSwQMJSApQBCVh59kKhGCD/4z6
l/GISSbnzqOLih9a32yDMZT/61fUStOXsSR/msHmk+yweFYhEAQuCNWXFg11rqHVGi226P6pFuwL
YaPOo69YYKLPF2/VFfEGlyfaPt6pDQAwZB7kPa9zHdUMW46/TXOAwiep5asXtQ8jxv/q1z+5nGWV
pERfyOpUD9GF9gvVK3dFYvsr3FWA2KBFmFYuNn3ujsURl6UvKO+9TkvnfJOECqbnwpUc8iVf1A/Q
3ZNK3Wm7xzAhmsOkuXtMRXr2n4lr4rvvcZ+CqV5FF7kT01XKQPFW+C5dGG1/yz/919fFa6Xbnz8u
EZzm1MJ+XbvZI5wEww+uXNfWEclCx3SjLprV7DvPB/VzpflhhH3uW5bkah2PkQhCqKaa5NO/wvk7
4AsXB5MAxz2suGcDDfo69/pvJNt/eK7jdr81YA37PwBI7oxf4uRXPuRcw6TiQbHcD1u/K50iI/CH
Gt3rSppa0uy2Lv8/UiDGXlKFUO4xUujY/SIe9vNxdbGAA2AsUf5H3/nx88DH/RdniRazYLTpIL6J
ZslnfMNlXQITuV1T/MgluiVi1Cyb9oLRxroOyjkDp5gkvDhWqDdbWf16Zs2pnsk41ZM0hyLDdhHS
VGU7t7jNBRiiCaEE9lx0FGJSZrkvcuEdwtO1elGvvIVULrYeNCHXmWEEMQOHoTELw8RAJSZ+ktmN
XLMfaELYFNKblgNUuumujjHjABC7SbDoczsEDiNiWTrtBkiGEbOKEiuwb8hY+qDLnFfHdVb8wTep
9g901S4Eu96tKbi59Ct6sZl/tM/v33jsipgbgSyb4HLw+WGCURzX5iP/5GTjUFZUZg8WV4eDjsLX
bXibdIBoO2ALmtygQ+nkSdYB8jbUl/15Efkp/zUpS/znTnDtykwR2Y15gGG1EiUJYQUoPSgh5mc/
4JMnA5wiG0LovBtWYQTwUXeZlXpTNKfJkiEFeXjRKUMjzHumu5JCY0ii39RgLTXGtMLk9RCMxwRW
D6jIA1HzCUpxDTYdiqDNRGWU/ECOIsFYYS89jk8sSOEP6/7furfOelrE
`protect end_protected
