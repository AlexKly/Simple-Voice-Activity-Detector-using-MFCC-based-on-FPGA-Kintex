`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hRIovrUsnBxBXUuLxVRS+mJ6gjQTWU5BgnftL7AlUpCi+oDsfKiA2dBlt20d8vRSmxzZq6htzycX
O325Y2lVAA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kBl9IdCIM3o3Ki+q2JZ5+BFjr679Xv+VcTquxmCaeCn32y3hfdQdmARjalK3OvJ0Yp+fFlA+rOlf
ia6zlEba7A8ixmZBOhvgpFy+epsIMarvXQk/DgDU2mlWi0tgSbBMHckaG7XEzdnYgK7yUgniJXbW
95iGCd1eHumcPV7nL8Y=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rMTI4EPuGy+XRyQvnouX+OUf9hPjA9cf7RYlXSDOSVku5bMEPyC4N4o7Odl7kwNYb80HsMgDd4EF
Lt7Zb/Z6WOSipNVP9Gf0I8gCz6hf4jNk/hVItZlgCHueVWrCemidbHTvrYBaQdzccA4qVXPYIXg7
v5AGiPv4AeHkWeBRF6Q=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wYI8P91BXQv8F7FCMW12ea5EiOrkEtcQMiYRgeKY2xTCszunB2zyrlpwrZw/Jt91uMSdzgqyXFUc
FA7eZPY46UU3bQzTowpkuDMY9TwMGOmoKABaPnO1l7W/PRnFyNHIYnSfZU/Esx2qoROUGW0HzovV
jM10c7eRuA/sYt8hQJpc+4tTX2qZkcLNJllFuN9nOknZ3pJcUnjqJf1UR69ySyUNH2ljDIa9KkVm
JTVkFeSQPNrFruhWOqVXNHOLvBLJocnrkykem+R+SyGEw6uEFlVR1HFygSlk8djVaXZlxZ4CVBkz
bS4Cix+XFQoP3HuIMDiwRskpb8Dz0hYMzV8rXA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XJs/oLDTJq4I7uFnRGdtD71df20/IhUx6yiZMT2TdyEIiQDiGwpZwBz59npVbSgvBrEN9aSwt1CT
3Tga3nsAm+OIsfMy7cfW9Wk9T5be5cYWmRUo0vuc6+QVHFh/lr9K3F0A7wHZALhdPR1XNLSPzH23
EGCBLdyconZUaIvucxBbnsnYbZWUnu0NGr01ljwIbuOjZNjkIhtMR69xxaC1YH4Tfrehq8gnxLw7
wM2mpqeyOkty1QxUzhT2VCuG4dEak6PW6PWGx30/odA6Drw95vNErfzUrqlQtEeDdm6Bw1YNr8k1
8iIw3u3x6UO7i63Ke33Nsw10TRNwcjCsHlwl0w==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ER2HyVPWy0Q/7TG8rQ8YfAgM47hJSBvwR1ElX/OsHwyVFv9BvfQrcZLpVRxdvxmGjm454/KHu59l
RA7LLZBzuSLwPvjJXqEMMnfuqTOWE8CoeO8160Oe898UJIIUt7jycJQzjxHmyUv+8vVQEWE3xRSm
xutQbXkb+FdMQsR0+1R/rP8YqIyjGO+DqWGmx/4WKP3r/yBQW0+cGBDSx7Q3w55VEnbOA3WMglc6
4MksecD/85SwcJRrdR5ILZnjLq8GTZUOLax6BSZKAirUsjoZeflBscgwr0GqE1VSxmXQwnaKeP4j
FrV46LgwtuGpgi2qmc1sMfMrj+ZAwAkAMJkMcA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 168544)
`protect data_block
sTFPVpGpXtoBd+cMsjynHc6zHU8sci4wuScSdQgZjrQh2xj4e2ogxM5/5JHDIQr++EJ/QlJ17LvM
GB+rNZqp8eQA1N9aBangdtlVnAeWD8Do8UxPYiB6JUHpP5DScpTXyNx3DquqXxyJN+QYPHMBR6ES
mbBCtrtZ3x7hffn9Qjbub3otYJJb6i9vfyaPI+YrYvhdQr+irILjo1f8YPLZTHLHhHXp2jtdmZXr
dvekxqUDIowMiYIJ8qNRJBjXTbEJN51oMjd7mboM1hW2nexe8thGdYTcUY5nPLn4r+VQ+84ScI5Z
WbcMH2WCiZjlMBOhAx4UgJVNMr9e509ArDlSXc8V5xI+SYHLGgZZulfnv53kZAktmHWfxqtn2Gl7
wTvm5muRrYtV6GKc2z6VaC/UuK96OQk5KXETwFihf2LjeqpfbfxtyVZtXaZ5oNtThSOOiH8HLWgJ
hNlIYJHHSZ+rxrxpBPpODVyIWBtp2klxcAplsWHVj3n4BuamlAm5gVGG6y04out/7hfhyu04ZSda
z+onLp/xWy7iiP36eWwbzW7S98VE0mbM37WV44ZhxzAY40Q4hTgiVbJHBFhztCor2QIiaOfN9A2s
BjxLH9vC/yMd+W0BHS30Hsag/GtINPMJdZVW8p1aLqY42CoTe3l3MihYFPuNQjs/+rkdcc1UB6qi
MvWL6lVHHfOs4eZ488EMlAFGJLFQEXR4meiNQ+YsUxEtlExjFCAiLSCfePf8ssl4aNnYGOXl/LQZ
mkxQhn2fxGVuk/23lXieOU5P8bgGV4MmSIlj6VdpegZ36d3PV6IuW9b93VzKM2rrNLhwJq2dgK3O
xpLYbz2ePHsk+YQZ7lv/JS220GXaGCZoYFkuQRBvdr7m+CxUPZ+piLmR2mAnoOwpykvKTxl3ntEY
bthsjVS2Cg0txfvnR+7JsV2n0LRtY7SRXJZQJuv+0ejybvdq2YR6kFV/c/SMvJJBExNO/mxDdz/M
GJDoTM+2+pnqdYGsbE3WUMfebqAciuIGXUbuMubB7ScRjJ4VnoX8/7rhSrnKI4hAyHScMJuIg2Ik
Ho40UKA8a5U0asIj2Kr8kfTitowui0SHHVE2GGRWsd5okKwOWfUOP7QDtZFAez7os1Iqf8MmkVuF
1YIt2H/z/Iml9NwERE3G6b7kBzQzQFbePw1hgchkrou0wRdxHhpUB1cQgsdOc/1uPi0odWW77YgO
zeJUaQvErZ0OgNpm85NGaNbjFZ4TphRyFsZnhM4EyAitbAIuhLN3+eldTCKb7I3/NGdjve1ZUsXZ
M4HNYFkqrOmMlu84Qlpvk4Ie7RVrsl5d3J4kZ/g3MscGOCf2E0Ei4JEj0jOfj7kp99yyjBvB5VO+
gXBNoOjQUBigNybRr9tYZboauusqQSRF/NYEsHiTmIn/Yp5lJ80Ycbc+2pJyFviyVDLIwVBV6fpN
amFLYeVxbPIXDkP0qNeXjNJywxUT5tUbkRqjCSp7xOlb1gAQYqb7raBPeiQJlH3lQG3IZOoKKEUj
s84YsSXjvbY8Jgl9BBPLxpvERyIIMVgDQDyBcS/+xMu0NYIAYx0JrXnnQDk93J9IpeSjfpUexyY2
S+OnW7BybDqHYBzQyZTBxq6gnsxhdWoK0zSh0rWx2sajxYNP82oWI3Nk9tTM4Aa2f/GaF7d0kDcV
btIIpanPT3q6F1crlxGFMzANi2js8CVp+wiuNDMdWDJiBH2KofIftgZ4p/uzqX4foWAgP6V6GEoD
vQf7UkCxULwo8VU6yt1+HZLDK6B1cNtWtg/zijwFFWSxLJY7aOFCCAE7w2q/Q5lFRXP30AzJnp0F
ieqI9v+GoBlVNY7DDyWIgk7LgGiF9nHKQ9+ZcATFK5pWpkGJXwcUjhgCyf9ou9Mh/PPGgouVFcbQ
Bzc9aLV2z9Dk196QfFSYO5dvsrUrE7XsTFZ41pzGuj8U5DBVhkHzk7gm706hv8eFWAY2OSzVYuOB
SJ0slGxprF2wGRtJUv/c+7/IFoejSYFtxYTDqOhcmXIGA1e03A58XGB7UvpujMBjTIUTuPMO4lPg
R+Bdky4btLQ2PNtiR/IbaEn/Np96sijp9q1nChT1CjUrb/gnJHn9FbVpa0k7XIFv68/dYj225VX+
gOlF+GRMBr9Dvb2ehxhM9gkSC8XT3RhBZ0afjSrZmKe1ME7Xs/4JFFA0hWT+dLWgE2G/Qz1mKEnP
INdugPMZpQ9DzCQgEJyFfLJuuqiCZ3O1boPpzeysg+wW7Fs9RAKRzKcWb5BTFl3S+X1pdKYpj7gr
3NckUzBO2uVkfYVULSTx6MKEYiroi5CYTXVi9k6FUv9u/ajekfko3rR7txxSb+lwr8fD9at6QKfX
mpgNAY0iTJxo5hfROH4sZIJipciyfbIRCZn3fahqujGCsAdLpA+kMw/Ry0D1NYz08veVJEenxL2H
nRcjRRoWFv94/gbZMDAHOSWz/icmnniqDdqjW9GGHvmgLmCeo3Sh7sgGtC//QD2YjF8hQTtruRW4
Vu1Fkr+eeQmy4X+RIf8cX43XGZOlUFgmzjwnkU/Qt/GGF1gd67+bzOkWcgKl7qatrdGVXNfC1rgp
TqkZMcczQgY/unhQjbw8R5wTomi5Ex0QERmny1i3iOGuLM6L9P8+ljCLtVSDpd7Eeq+sUxupq0V+
r9EK9db1Aldls6DD4vaNSyr8ayjOuIVeIhk1pIO3hvu4NsLLabbNFcQ0IEdmoHAKYeCqoXJ0Xmo/
9cXgAFQ4Ah6/O10qbfoBBoE0AMKcCjIQjFEymmdF/VB7ajsCKzi8T8PX/GB1vZzoeQDVkg4MoCE4
Ce2oqY0uuwNncDf4cbKIrWue06EHFOZBEimSchIX805I7qDl1K7eJdpKj6QxueqjFu2De9/kQ5er
XNJRBdhpsghvk6fj7FiLIHQdSN/4KeDMyIYguTPJlPPqIcVDogYXxEUjYh3ujv8sEGAlkvYGjRhc
BnJQ/JW0cD3etvQZQ+zgDOMv2YwXztpkkEMIPNDQPSsgQ7Jktbfe368ewlyNwAVPirB3uhMpBNNR
8zQPAzBYfyH4Pw83vmi3lqT1rwvnrmH0E7dK2OBoms0MU8MUbF8HvYdoM0I2GX3Cbe6hQa5jfbcR
BkCnmUOibsBC4xJ8DF2svJ7tFt/HcsvlUs1eV2kl0QjP6u2dmibpq65DIkLfdYJbW9L1uQuW+8zT
O2VwOMHVCisgw31VF0htST4GxXWQPwfqlzKjxshSRLWf0yp+aaGRj9j22nVAtjh1Ugfgd3YNu4/w
8a1A3NK3cU+cSAGIbBL7Ps2xpVnEY1uj/EOApFaQ+8vpGyZEXoVJvelYGMdz1wN8QPXeXBZWyBFg
cpvRngCzCB+IW1hLgEjGpNth9HA2WYFel8mm9BBvMPyvhKXdgHupzHMlxA7xTpl2xO5aUIX7TyRx
jlmDM60IuaQNOvS4oWNRPZ6lWML92jneSYynPTSRSs47P2xjL5C3tUgelZip66knml3whaBaUbql
rtZELKsVKBZl59b0hTldCrL6iMnNgipnaPCvgeP5XRj5nQSqIOSDfVMFL//tbBoj2ZAcVCpGMQyf
UybUBKlxMFuosJ8OWsI/6PctFjM4hnYIpKhWfgUrBgUI07YQnZMxiK4sXNP/Nzxz7qXPB9brzZB1
vlwotWLa2OaV142lIs+1Pfk6H8l1ThNvTgSeZYki1BDUGqT8x6Y/4h8sU2R2Pv2TfseJdtveA/RT
VZfyTC/6UesQs0tTemBgRuEG23jI6Q0PYfCL+4ev2qob1Y1WW+YckL1PQvxP6vBzsR1yvAknLqkN
oWa+ke9VTNshp+2PjWexI5ZIjDA9gCYugfvBCYDTOb95oe1Z6KpnRX+wZ5gjpbx0fMfwSM0HolVC
zwRSZEiF27bvNv769Zmscbc6R4mDO1+k/PJzKyGrqHG++o8QPWURUkKIk/T65kW7rnyDsy8e/Q8s
bbrZ2O8XJtkzfeKXmm/XdybjiT0OC90qhCbfLMJr1XCXSWbSgl87GJMr8CDqwgNHvtq6g7EF62DA
itTqKxIQcg+mNy/wmfA5JEnYzMz9YuBjIbAegrgKG/S7GaaJu6fu+Lvyn3qHMQrYAF8KCQDlPxRJ
gXwOUxStItrm+gCNiGfJFXO2kiiSS+4lT9e/D1d/D1QMQyPdSWPJTb46CuA6VHmguqTsbhwx9bgK
aVwxdERLD7FctYaQTNZT+5f6reg4++UY7duJhOXnRT5xXQF4jyOlR+n5jAujkHoAa/8IRuSHOakQ
IwyoJPjPO6YzVQtWs02Ptdz3DrIpxxiGHi16tpimfDxYZTUD7Dt/ssI0WFu5bilZAt9i2zK76MmO
36kj6AaCMyOLBEGB8xBWD/0dFGNvxeQpMUWgOm8LwSIZKBaNt8VhloMEEbAai2LOLErQ+ZETAdzl
jV+uZNv6+MfUol9Fasj+6ErPub7eeZdo4thTG0oNgd35tefpKjlfwqJx0bseDTUs1hUllEOoM2eH
lydR14VAueWi51K1XwyUhqjLw1bN7vTSr+4576OvpZ+K+/bWYptpAqbrMp9lxWEVWIwkPNY7B6WT
FmsK58Z4s9rqt5AdjImTmbcnkE79vZiOeMxYUPggVOaQ7lxjOmxEGZz2SebAZD+7s4MXoxp4eV/3
PQAvzfMHAn8HdGvVQvYbGLTDupyv6DAfZsCJBFC/hv72CHLt65x9IUORZoHnWvE+me12h/x8/kal
0mZWv09n1GQCubs2MtOTJoWoGuX5faX1JLQ7zVMoJ8RBgb7XxBQjFT0RPiR1JXbGk1Q9b48FTszR
rlQtHYaqx+ArF4ZQMc75gHOE4OYeeYFlEmUFJ0yGN0wARq4tcoSOjlr1sGrg3aoBP79/L7w3zWJE
TKhA5La5ImrQBAkSP7dt8hVq8cE+r2fvxs+PAfhea8d/+zpRSyBCU11HQ2k1LH7cDd5tTL6mT3Hn
dc1NCppqZZCgaW1HcwrsrWOTeGrOBtQQYLNA3rCM1n/3DyfUtE4c5lpEKXJehnuKUf00Jz8Es5mR
p6i+vrUYoUBDTNYmPxS7u1wSTryP/HcIYX+6UB0ePYUJ3GFnPFWS032nLaXPPmshEaBX0kmtoGqq
l/nTQFPsPLg4qusGvRKpeNRwzFE4Pdvz5VEp/KIHkBhvCwY9zYbtp487doIraq8fEr1qh4vobQyo
Ns3hTwCFlUvOWNIq2xa4RkFCVWz5QzPsrsEfMFURLG7TKIcwjR6XOvRjE/amdSHetABFmiYzdcdS
D4OFsreqmO82+8paojIOQs/Dsd0ENpt2LwWIjNIbgjlM9plB48MPOEG/0tP1MPqqNBv0Mc8a2hhH
UAsOULyEaQKzL5p8jtpUQtoFdONqJeo/2OfdHoyLalsGaqvqn3CE8sICJ9m4mAHAwzjt0mxGBsvN
F8NcWqm20jbVORR4L3VfvzuNgFkLBggG7zq4ehn3b0xAkcUomz1yot6PrlDDePNTlixqyFx+Bmdt
CrjBomxsb9OSMKS7QAklBEoAw2kZmTGpSp+cRSXIHs2QG0y8qxvnpVjPHel55czwTiu9hbORm5yV
z6i3HZlshiBFBn/hfHYVkuUhYgyMG1rN57L9UOvhrSHxAgcEZidz5sF/5CrreWwkT8UMCNJmksDV
FB/1SfelDMDW7JlrV2dfil8R1e/Arm7LJiV/5r8dbTwdmVJn8kKIpxTW4pJgwQtZFtRo76EN0DlE
ogP7h4yUFza4QFTh2CwVXU0YP8mEbdpSiwtKvKWqH6txJHtaCRBirekUT01hF/oj+z1Bb8as1fCz
IExm5Xk9ixiUVaoc/TTHFmJQIIEkNGGRALv/53fb1BWBiG4SKqzj6hXlAsql9KdrGu0yLFElH5oH
lJNElE4Vu+1FZINjgf2s+NLieVusFrFtOv3lyKl12FMfPx44GQQ+ouOil0Z/8DFtuKQKHccoiIMp
9ckzZhmIEtAJoPB+FC3I1pnCPFnCGvuMg8Iqsb9szM3tOta0qRDXLbtz1KmvI6AVVfL94dHFBIke
4h6NxmErXQvBAuzovqFpvWhCcHMa+vzh/YaInK+dr9KgxSKXuKTMaGhm0YjyoZ3N40QuDAnI9kt0
06iWEY5+Th/9fWz3kL8JDbcnDokjyVLHUaoput6iRg9OcAXh1lU5ww6BjO41TFmj2WHSYMoCFILM
P+p48ZXgIuNMzwYqdVHW9sVDRQ6CYNb4EL2X6o0ls8LwgTCOj9nGZpfIpH20018j0kyshqRAktT7
5Z6sVVy80GBVEwl1svIUCwvGdpKjuNqL9JuJxHw5ZBXHs9KjP8TIFPQwvjjnU7LdqxWhO6qgKQL0
NgQF5cBDAZ4elaGC5VJBekbv94oUemwOKWkLMxbw4X1DPOprAVdnIjrtrPZFZJG1xw8nkJvn3ZoK
+SwAde4kwGDe7a02rJ7ly6rYgW+7fEnILA2kjyizYvHz/1PypsMnXnWdRlml3ThBjlM/zzhoIAa1
ETzGBfK7i6icRUJiF7tdByaPx6dKN/+I+OI/ePpoG85Dj+5k6+RqWyaaZVUjZjRazyM7iYA9F6ya
zz2qNNlPrVAgQPSqB9RMYzg9HZc9qpqIsTTSbGCVZOEiPM3ry+FkWjdSKLATe9bz4AtavGx34AY7
ln8Rsguwa0FS6vUaJjxvNFq1XuCWhSmAaGInCU3cwTdaORwuqX117XAr+UZk23LOgV1tAN26IPgh
CX/vizGufLWnV3b6jfResZ5Lf0TTKfYz0Q2EdNBTX6g3K2Z6zmDuovtbc3w/tNfNia+ki0po8Jjg
ssq+QJ5fCd/DxnIE+RT/j+FBs7ZXt1JFesS1YyaLG5B+prmdBLkPr2dGm61knoj0JBdv6LDjnBAn
8YaTTqQJuuMAXhZ6ExBVstNFjr8H0msvR7socqN6R9aavhJiiPxtBu846VLDg4D5JUql6xWOYMwQ
nk+ALTDusgKjvUlM8G4DRhDXjnn2Nxo+G56yXbrpPaP3c2iIst6sJPAfNnwrih9JtryP62oe9WHZ
lClW2zA/BlTqryORlq94lCEI1y/3UYzeONvFKvgBv5O90+FBJa010XG6K4RG5GPinXV/1g7aMmlG
2MAXAXnSmeSbZTj+bilGIvssuzSkIumLEraIeBfpL5N5EcJUDW+L82JVW6gF6kMkTgnGfg8hnzS+
MgKqnJ7Ux0tUUDHlDe5ZtmdO5ckjJztTPNrilDr2BVOL1LBRgEdMClW/6RV/bzlmJR7fs31JWhT0
Kok9QZ+0e+2FtMoa9G451sNKLdA/1uL2mTHjx4smzgTGaUk9K9o3dqT5ht4bqcy8mRC1/JX1hbW4
mQKSmzFWkfc7dq0HxnIG420QJDzg9xE28ddT10sFTpzOyOaGygShS/BYZAzlFzyg/EKo43MwQnwr
UFA28HNDEjRB9kdrHAym/VRRQ9DVIT55N6oLZbJo6m6AbDQNLPGE0OymqAQFNib03KofUJpVVAA/
ZFBlzLYLi1wm7ku4k8MxNZglrMlXTe4Cd76Za++z6ANaEbI/jkwS9YpOyHxdl/Oh+vMOG/zDzCZh
fP4LvsoREj/4FVujNzwdQCw7uxm9G6otfJhiPVRqQkowNT0CRX+Ik5AG5NV8Nv1fIj48yXZc9Wyl
sEmGvkh9g/r1FxTr1eJ57V3qaO0uqg9jPgJIQXBItI+lQvEgbCrvjXFRGMa54DbYWr2m+W7dz3qn
gcvCO1hREQKYmwEKIUhSyqj2g4zyTy0pKUQpvmijSK/WPQXBTiyDzvVul3pX3OCgpIR7PyxmpNqB
8IqJUiUwf84wofAHvWqnuBmr7N5U5cQVzBPygQ4C3zWbG/vxTth0x0eB1m6SqYwEa//PZXmAiGAH
eTT8jMgMkZfc9JxZJxubM+NByk90VGwQuKR5otPgrc9dhQuuYcCRXowRK/DsqHE2gE9ryNLn2qS4
TTz5ZwoQOxVOdktXyoOwr6l1flRT8p/hK/gLcvXW9DaBnRr6SRS5ANaP3VR0DKk97SQT21bg+SHj
sKvZ0uEO+duSryJMvI0qgoetIuXvAAM6CCzwSO11hhcdr9HXLnwwCP+/o53jofWBTbeMQhW//Ap9
WkvwTkrJsjTaEOCkCvHrFaHUOwLOEYBsAhczq+x7TEB6NKMi/E58naRgmsTgOihQbB1+mYqGoYPS
WJEYk0RE10jbjZO4eMdFK6GgVc44IXWFd0VXy9+5geEPEqc5gEnzZsnfsZ3ghyHhGcuw90p3SXy5
hjvgVzxLdMJrUDf7qWoYybScdQnS6412frRWzQTGMwiprWBpG9AawFSHc552YTDZloCZq3zfsPYf
JgB1iV0RANptiQ1msp1ycn3WWCEILF43f3fgKiMFniBAxe3wRGyk1qEKtxiau6aTE1gDk2q2+pav
NYd4IGpW4DQI9OBLpYKLPEsLrAX9PJK5UiwUUxvOlSAzpmmtpVOFJjTwOMaUShK4w4edwze1WjRu
u4UC9FFFQlfA4jADtzbI48iuUj1sebdKvNfGvbRlunBl+mfacPgx6QvhIh/XM4eksfcqYp0VxeXS
Iakso62P2MdPKY5piXAed30+Hm7dypJm0fsF3T2DW0/HBSYmWUw+Jrl157QSgdNNoJW//+uaRg1J
/sPxkGd30RYCLEyhEQssuVI2QjJFfJaJa5SjOXJ5WlHczi9+B4Otzt9FdDatWJigOHI4JK4cgLOW
d+AwVQR0ezw4GeUXVLq4uCiX/KSZnf61aytVavG7NMYHor9VDQDaZMq68xNjOxtSeBQWA4zK4d/d
o4Kh0c0Fi1CqwJG/hxrfn/ir4HG/XmqgNJ4til7nUzPcmfPoLdSfVH1p21KiK8ZLgvkuukv1BLRY
h/dY8VpY2mZ1OYOdzLz9MdMhra5xn6ugf6wK4VZN/hkk0HVJxKptYsPskdjLTrufWWy9/hgnRIg8
sH8ZFRaBoCMAYX6jkMH7uI4aWHPXHK2p2r8UE/zkXHD9OwpxqwKWlq5YMlGEUQRIhPWJioZXVZmG
ng0MFXCXW8BqasfeB7kS1OyuDjuSQl6l3hVrxjO469vq37nMiGqnp1eBH10ktKyC7uzNpzT/pxAh
A3n+Xyd//VwxCeSb0uao0ICLl+MqSEyBMAN85CPdWXnaRUaQOdfKT+6DPSXzulHAmUU3FWTpXIaS
hsbk3vlHfEKwx1QJjXkpFtZ+45AGPU4aKv3cVUmgU0fCW095LYmXeromkOtJ6E9kImtl/a/e3kfy
ACyixykqnbJSlBOVOAqRTQ9PEn/GsxPKPGGyjWtS3sahKGxIv7xNV5DxKFVVCIzglZbELVyyNer2
OP1HzjK3iv5mOKRtzc/wBMOsy//B4IQiFWPiAF31250NUslvcz7qCPiuGsrLEgoQa+87UockvbFj
FWwiZauBmRj5BoTOIUEDu2NDgak+15p4TyJM6dyR9GYpmovVnRQ2spMwXtLoygyrr/qAZPCtDkFn
yYBB4Zx2pHUYXHrRw9O7OVGgzOM6VexSt2PxZY/qXUx4YeB/Cs8fh/nCWKkGtVmqzQUsr4/Yn53e
P/hwb2aPDumIClz0h/ZSqr9F8KeV8jOdLp+BrYBhlkP8y8k0NACRYk0fs0jQeTyG11zkEC9me13R
FWsOn+qgbYBdOxoViYclA3HNp2fTrYCJRhz64H0iHEQpHJxK0oCK+qZOHrZgYI6phHzgYMMhPp2C
EkMYSrCd7iI/4vu2+i5hTl6EfsLWOuKrKKHb8m1N8ofrr3K+z/vwR2srRl4PrLjezH6pBzJRVAGl
gn3FnW0WOh5WUU4d2vx7yGd+bYSWTi7z2O4n594adMXsUW1lHT4l5JMQnj3G1E/RLQCTFrgvM7ek
VN9mOozURSLloAINX/oUDUaFnHiB0qb1qqzZVCXkT4yAZkWP/2JaMiaheMD5nv7mt/Euv8ojGOPQ
EP+RKiq7r6Js4zIym2dChER7a+AgdmHK8DDD1PZTFix041rJ3c8K6ES/zpTvGBJyTeZV+8qmhCu+
5Rxr3Q8qA8VIQzZ3pvUiTx03W4GE2LSg8GruNPI+ZuEcSu5yv4Nvj4IALx9CsTN2Id6Wq+JrLCeK
HVl+uxsTiKYhryeQFVYE0tODUmsjDvJ0YKhtDLFzlYDtN1t1qVEsyCa9evzlH1ZCL6Kz9GTmFuHb
Vtb/6OU/jlU486n9FvLBQRmFhAZGezf5oQEHwCzRQQ2lFR3tX1flIzM7St5WEk2O+r5chVk0EeZC
MqETbDx9UhFJ+4/6igt7828GWbWqac5FduLDPxw38C/Vze4BiGodqhexUW2ssqgL/nituYo3eCib
yBKodmyzUW/tWOc+S8Zb0vqXi7ebT3gL+n7pwSUzyOjldbSfXrGekh/iMq16T/a/mOh6q+Yx3cCK
xGXYUVMVMxeYfqjsjMcRviM2F3e0xhwkwNvrVid9ZdXk124ckRaFj/LNLKb0FFX6p8ozY0z2Ot7Z
xsvKLA1EPxDiq21/iNGeOI1/LdypjLC35oWcUv62y0dxsrP9xwQ3jmzfQZK2vHd0MYw8ahrzvbh+
OVJUhqjfx2AtCxjQbD5VMtM132OcesGVwCCORWmtoz+rGGorYhXcTwjF5xz07Ly6SKveOm23Oc23
XFcjij7AP4skq+SmB20Q/GOcUldGp7sOMhnWEfKCYMmPUY5YCxzpDGXbUEuKz9BJBdpLKXH6E0AD
gQyqIPqID4ic5eLkBUyTBYLLbdlFneYKkD95QKBxqXmrkHZ30Hxo5CtLKKD6U+izKyVKu9V7pnwh
mw9O8z/85fGEYLz4d6SwaJVplPseD+xKZ1NtDMirv+Rla/wiJKiKm8WDoY+/PwbRgx2grqphj2e5
n9N6PwVgigHHHavOsP5ROa0QrsXRHZXBKsEUx01f62onzW47X+6l1BS839KhpUnx0Fa+Z7BNpHT6
V8+vQccxiP8AIDHn+d49dgzHuU4BQS/pGMqBXz8LfA2x7YyIEcdqu8pXFrcdCAoEVOiFtAGsCVuN
ZNyZz0MiQGVjQrNb+KzUnd+RYfs0df4BvzqNwi6GFF1p9CO3MWm0KzmsQs9aqa19BKGJayGlJtmu
y1kfegbqUuEavcV0OEDxVQ8MSTyB2WZto/JrMq/6Yvj0l5vOOHcuSOWD91AhDoFiBkiKViKvzqoz
Zj4fd2BFcddtGlM1RtOPXIfbBnYDcH8l6+unr46D3XsGOtbsUJjFafTHnt3hmbY7zDWEiskvpsOW
TW+Qckwzs/Kq+GiHhmVFLh9YvhqPOmPXk/P6XMH1irsgN4Jxyslu0x0SBEqn6Br3M7YudEKTf8Lz
s2BcexXiZcLAoyYRv94/oZODB0+xz0Qvzr3TBF1vAEwoKPsbDFTZPEkTq7spitQQaQe3KPaHlux8
Q1/xfEgyyEfnnF2md+3/9rcsGddVQ5we3Dgbczw/F/l5+6mvXuMUXHs4koMM/eNQVNIbhgK9MFfX
yEC6TZAEzuIMCytmrG2iltP2TZpA745vaytGrFW9vi2VbkqDy/QWyOSAu0IsMltV9uznyQbRaZGp
AU3FiC/2NvfAjCsrde/B7UBC2nYcGmd9/2ZGvjUWwlJPCysY0N1GBDiBp/wAbYqbxSTWxWUtif5e
pl8UB5QIUCiHucIWhdOfmm/iufOrITzq0x8eiVeFqeA/EhuPbcrfCYd7IvgdF3yRYFtdnrHA2llK
7LuDmgMfGCu0n9m8EBLkFMfk6bpGdxUc0Wjvy3BPeH/dO89CatuW/BrCP6VYQOgtsA+m9FVTgRRX
XRk4tr2ctDbXFn6jsXYsoW/3MRgNvnpxCGmtVRhvL5dkGqft99SqeCqd0r4gt9+N/K/Odn3KRDL3
0mUu9UFhhuyTvFDxfcW+X0FZYFo12HtDwiXguOlZPYMcR/u46ObCk/U462uzAvLg6w90mLvOL054
g0LD3Z5GAmtPWr3yAhCMg0qTb1AtG5ndYFHu/NEZ2izJTx/ThygL+eJ9lIjEZvFk8irsENcxqUAy
hAh4b+9meFXevhO+i1yUy30CpWTgIXlfWofHcYOYOuX85jFcDBdztSR6KXNt7XoxMmW98052aA4a
L8i1H8MAbGXoAA6mTiuJ4DjMWzDDdGcVFoBz1wOAvvGWXnImyweWLIb+25Qd/0tgb3tKXVRMJmS0
EVv1m4o29Gv2XY7B/sG8EVYbhQpnutqwAGDXoupYaiwwCuLTgkggZuCzX2u0nq9Ab+WObeMGz7MT
GPHG8t+NLO0kq2P6CCiaPBIO2d3FwnsnVrHtOfo/ZWMPXcewyZfIIiEZZrfzbBbIQZGSglgI2/oJ
q/EvrC8uePSJZUalCOgJyxnu1i2D8A/hBTDtnF8P/71qJP61FBnoeIXrneN6RgDhnYnViF0C49j/
7C+JP1z7/nu9pvRe7qmpecd66UxDNGY+B1TG8Q4jCenVzySQEyQJM0N/4i7YI2nlOimBWjI+mA5j
OrM5SOD7UnpLhLzQn9/oo0oeiPB4S5Ucu715r9kl31jFK0+PiT8u/jbv7eePwuBO7qR5bP5IMRQ0
QR+dyYRBSoN6bWMSuQJL04jra4FHyR/WK7kxKvwvhQwUxkIpjGLjjHRYaIWcFNJRqyfbM9BrcdZd
wx68Pdv46HuDHkFVTC5As5EzC1YcyYdZQERa8nVdoK9E6dXS/iCbFS5g8fZrNcuPCQQ9hEAmP1ZI
Cd+BuuNWKj6A3HiW73vfSwuZ/ArsVYo/xSooFPkGFB0haK5z1dAkQm1qfPo9uNjIDGtQC9fHjJNM
iu2GZ0eDKpY/DaEwnZMPSbNo9/zzAk+3FpDL8gUAtEnhW7BIQiHPMGsmmZx9PyaIEQRVShT8RLnP
07LLSgo9WnsZ0SIlNykUoAiCnQX3rjsGqhvcWbEbc/ivsKrrmoeDoiTGpwE4DikaSOuKp6xh6Esb
pVI1sFL7DmfDdIlIYikrr6K4pTBBd9r9L/Sbd1a1wj+DPmWShbbg5/WeJWNQTcJmfs5MpYwH40/H
dYiIjVZoxYK+dc9DaQepc/C71t/xD66P6JJD07YIcXNnk3LZxBGpDkJptNBifzFJOrIgJkIKe9ct
WytkQiB47+zi607n2nvtEPbd6ELuF6QvZCdhwgmDObH/Y9hLKMhYMShssV76j1+QfaiANwvZDx2P
N9cmDjQ0M1qrgkEHLMf7b5gRYSpZX7EXpliNTERZwYDk15ex5iJI75Aq4tjjWp3NtLVh4MXhSMJF
Y2LEBFeQtTjEaerN8QzOqAwE7/mdIkGQX0mdLKezkBPCSGEd87Wtsp/sy6vJ8F9yWWAHAqC/Swm8
d1zJ7krIgwz2QscYHCwjI49P+mpXneVAojZg3wmiYZfAk+6/HNMIFPz+xLUxPAPuu9LQjUH44TzL
gucVf2uiXX1RSZXECIdbsc7AktdnrJRU+WiAZixdP//V09OuLj/rKycPqharaKDoIH9G0bXUw+So
xH+qkDVKNRHI7kaetfcdTAz/ys6/85nDgMRuxTlvz7+BpDPaEZo/l11HCV/QhW4SxprR/t9v+dFS
FIXMgwAuNsUOnY2LquDICntJXPEygVntSbTgXgM5IE3JVKBbtkZcUIzThYs7Bm8NQ/q/Pqrljqf1
18Ma08Z7ZVoS7SjMGbrRujL6Ne4or+sL5sHAuj/DdYefYq16pmmcxXPXdthswK/5Cw7Gyku79erw
7Q9gJKUfovqkHT+3QGs+v7o01/M/sGUuPMnYXq4eU/fIhwDPCzWppK5a9j20S621J0XCFphIlpsL
y38e5FNTedYHgbmC6eLIrQllroFw+VNANp3O0VYAR8EsFdwBiZMLrvTvARYu2Rb1vkDuZY6GNIeU
kyXpf3ZCJXYq00XW/UXldfSeHdkGtdMrloQpAvdRmM+hSnyuPQuUyxqAOMrenm+BbhM1ncxmiLu4
/rYz1VqP8wZml6UJeWKi6ueBD5sahMXM0SMJGTpA56LMeDnNeOelCmMlmRxY3Dx8iT/gx6XH9WA4
5UWI4hShCkou820W8x+2k6hnSv/hKSHWO8Pb1P8hFqJJiCnlYJW/g9vm8cm3tNiIpp9kZXcEJVRP
DA6Bk2KzA1ZGFG7q/luZL9FMrregVWfPyw1SnKbrwJq2VYhHFz2gvPeuI0tqE0mHZMbWX4L9nYMn
mRShZmnAo4iM9xafIH3TixWgkNILta1WrNF+SWnIN6m7dRo4i5W7mm2P21nj17jbCEsU3vv7aiRg
S7RAHzJhVst1DUAOK1bwgNnVUJ9DWYnKYToQ5mAsoIeKv8j2n7Oj2gTNVgAUm9lGGrnKup3jFYaR
p5Gf0328DiUtq4qJPue5an/iNRk8QUhrWJsD1pIN6JUgEjueZjL2JlpYHrbjrz+DdhLqXUFvlI5A
CqbsdyK+DuJw7xOHr4lLMzXTo3isekMwGXPIg4y/wpnOc7/dlDA+/pXBBQvHoNn+4XZbudPe1vn8
utoqav+vrH7BII+2U2lXZIpy5TVIxrYTRj+DhS5qGnh4WYNPPEqEdZZoGQPMziOMxOw8sNA207Wa
vQ2eOIoPXpNVXuiDs/AApBHeam3ERCMM6hfu26RXnk7KTITILJajhd535iYtwlKxUY0IWhBNDH3M
aWD7ARTjBMcC/AzJzjNGgAMRYGcjeQaXX1stNrD9qNJXlJzGGoBBZEOUG2DrWRFvw6w22RGgh57+
Dd+92lAiHKPXtroiNrQXHfh55l6ZiJrwAez+T5sAacOffPAWl8nqe3uqq5WxTd1COWtbHNZKmq6c
gsaBuf3tnPjhO29/C5UrM7P9Xw6cm2XGFCNEmRitYNAvJqspykH5LvoNPcttMYj1G2N5W1paIcpv
58KnPI4no+znXOwQ6MJ2WTahzABMFxD766sE5z9wXA5TskE/YNaq2z4pTJ7M4EbsG0WSUoFEWzpf
qjttu1eQQDFRtdiDA7CQhDlqc7FuU5rJWglAJf1Q+liEd3JMaEN60H1XWxFysU95OZ1iOVbiizOs
JctiSEi3wcatHekOVjoRftJNTMMly6+XSrd2xzUxZNHUZhwZrDDVUz46S3BFlifxKzZtJ+g/5KSf
+EhWnTyiGBCa3GOgoX8b2gDvuttNtvjYctKxpHcW1z7NBiBhxGDpx97AG88nksSKr56DEC1bl3BY
Ca3IHs1eBD00arOkqxjMB6ObN1mQG/gVI94e1yJA/mDIbgCoTaBH4cnJY5RFMFF3IlXkGTnKtr0o
77vsElcpNMiYq+J27aIwNEuQHuK5ACg2JF1j46mG4bC27Fxhp+biEjTHV9MGI/X01attmNDFkpuR
l8SEdmrHNq30z/NQblwZnVV/XeCesn6082xtPrjrsUpIVnrGEDrXkDRS88QjRrHtk2KEf2Tgw4L2
ivOWQZk95hHKhHmGcbH5yOmxelfDkfsRHxb7y8oHQLEkOXqd0mML2rdAfczjS75ga1dsA9pjLyE3
BT+HeMzU1kSpRlDTYo//oKl8SDYzDFwiFwopWpI0r+rVorD/1qjq3lbgre+hMAvfgkQ2fR2IJKjE
HZY73v0inDw54wq0vXyZgHhVc40U+0qIEG0cSTelU/3ERSDiv5dliRMh+oGVHpbuueXz0d24SLkv
UJD22O6OEO/S8w8uIHACD2N1kupKAmNxxSeodtA164mcgeRvJpRS+HWe7dWJ7GxNXBN4Krb0fBW9
MfeYwLCKdRBZYChZmimfKyt0cLXoOXKefYqQoWZkl3sDE7whu3w98aXB8ksz1u9vwwCf4/vQYd+7
GYGFEVp4UMWAc31WHVxY0SefnSIZFI2RrXv7JacNoGzBvJrydR5wnP7kauVYjgwlNymXovY89aAp
t/1mABwM6NBSGQLW1elgSBimoTIueqYGtM6RYyyY1foCWKcPzcLQS6My9Utz83gSHVUxSpjh3gZL
MU0KrdKlR6ErkQ25QUnCxJkVvztEjk5TB4OlZnTCyVZwI4qYkWY4PhnCn3jbNC+GgF7h4AClGT6m
OnLhhTSJ0xJ+WrzD4Udr5BuJUgNLEpIeqzuD4cnFV/bHLCdAHAN++AyL7tUFQ9hP13iraGAPhqk+
9oxsmZ/A6Kt5qpbU6AqddcP+gQYH2XprcuVL4bkq/0xl18DJNtTb8WZYXDaD9PAerRGBiiI/FG/o
+n/Q7kY0jA06FoAXfXjolyO7BEwgBC7rwxbV5PZAoHtRMjy/7x9xLnQvImpysCnWiOABtw+V+yPW
WrHXCWYtJrOHPs8vZeTqCzXVHKqMhfesC5yl2GcuY8X5gigo4LsyAVymq+KjL0UYl6D8QGOe/LKW
ly4SYSds8Iy84YXa9qnwxLaVmCfx4tgWiDgAlXqU6DD0GcyRVao9wXqcoDuZ8Jp7GqhJ+ZaaqxbH
NCmLgHIN2y4pSnjvkT/TL7jezv6N2q17uBioxwKRz8eb4O69MYO6jq1veG7r0qc6Rg8jXIWQkZlg
aDfjgzDa5F/YxYK5b9dJ5qzg+TiLS48jaO9WG+L+6PoTvohcN0Sm4/ZomxQ5gSHLoz5auw7oVtCb
bF+Q6D0GM4QrL0N7f5QPQEdeNqZyre7gfD9B8qbpL8Dyb5lLtgYw+sMoW451Oy5191BliqZzm69U
rMTw9BMVIQHFM7/wiogsSBDa+OhfiZ98iS4qFywKs0tIRL3asqvuYQacPh94ngeneJOHJd0egh+v
A0GsFAM9g4H6JL5mbmEyyq4GI1JO8C/+Kwiyr+eRLp9pmug3iu+5iMbg2U3k3Jnlb0DxFmmSIYCQ
bUuSbeKiikWP0mbd/9pe8nOVQMgwaKsmhCurRbNdImQV88z5QZNVgSNbc2x74M4axpTvhV8wZak9
CIxNccqf7d9hMcq8mdBg/v6HEieE5Acpj66W9UGB7zpVbrFpIaosLlHz6YMTylatkcesgEqKeqiF
8pcimftC6PJnzkp2Ls3vjaghutQja/5pbQW8T1gym5++/VjmQ/hir9HruTzG36nnoYz0p9F9HJLu
epmHScrEi4PyWxeMyaG3VC40zRpaRT+HEMO6DhWtWOGdoXiOMFYDtOq3xpgps5Ar1tdRYAX82dvT
l3J3GSsjsbTfd7EdL4FeNj4F13hKybxDOOXCmO57olmGnoeeW12/jMMbJFy7RKb/2Tioem70XhI2
ndjQ/MRp0yx3iB1GK6rIgJL7gAEGSBBqrCu+IhDa/+Lc+1j75xrEAxo1MYppHoXyW+BqyJD2XoZQ
pe6LjtBsgt7oqilDBFZEIFPfFnIeGWhBfUD96zxoKVWLIp6RERliZMUQFquNdIYFsPsDfJaPKXCZ
yTe3nIytK4GK0XCRDBLvc5XYnEH+3PVzQ+jkL535R5Sx2+0fAbi/kT+94mY79xrPF5cmWMJ3nWFp
jMUH0HE/5uoGCD7jnhZKgH6LzBWRjU1ddXnMZbKULXO4ou4HjRmZf+yUAs3IB6WmGHHfrPoaTg9g
d/ZZcQHtUe8QjbhHkbapsV2PK/cGMlHuQpDW69j8Vqspa+sVCSsZbCyza5tu75Sy0bjW0FqTPBRz
UY4c9bDq+YHnhTC1pYq9i40doLAU/V0rw3YeXeBoMY8c+X2dptqf+wQ9VHLoKion9tVPj4/1TuNX
RFh5H9uUqAgrEDrTFl5ZSxpzs8AmVH81oBYmFndclpyxBJAO/2TiQ5Kg+et9clIvRwZsRW5HWVcc
mezivdg07QaIWkJpWlgoBBCJoHTBc7h0jFIkzHWAxWk90ZrnPzG8mHZoNagYFMYzsngMt4yAk2E6
84bU3LVhuxy+wp1ukKf5+1VPFPVGc2utjH6aiZxXqqEIl8i6H6bhW40WeW6D7n1wsrFzFrjdMIS2
Bo6eSAfADjcie9RxS5dnnaxHpZwvuFaP7S6vwaP/hTIG5cSZgBwZeqwsY/aYopxO5ns26WAd7fbR
nxUICZLBAAVlhHQSHKODLBVgWNk/0SJt3CGRHLYMjXaA/5N8uNoKiRgiI9GF648gpg79Pzuh/IZ/
bqVUYuCgLW7duWxdOZi6TxvBsGCHTWV/QkvyP//rBd4EabswZgxfa7oahKqAOI+JtQo26jBCxWTW
Bc0pIN76fyB/O16Zpwo0RV6ptOUJPYDaJ1nQnUvx8dBYENIS9dDrLWd4JIh7uoFUH6Gd+nMxETe/
Ss7NLRRdeRisN1NdwzA0/PQ5+zM7qdQWg7SyVFLjk47Q7whQB+oJN/6VwEDN019vet39bAczOBCW
Hk+eM+xFACoSf4RT+8+cMS3UT7ThhqtSLig1iCZY7IsC220neYIpbSkISoMh8cnfvJpuMOcC/Vs5
+2gYA1hdR5JMVwASGPsNYggbF6tw2DgrXjgyfBRsOBlU2AWIFJVNGiPf5TQNxYrYKUQAf/w1BlFJ
xYab6eoiqWM43McflBYVJ6Achjhw/mpIYLfTKkBggfSBJ/2CeIB4bTtrgGvjNBbv+bDTl7IJF0aW
m3X20zfMTsg6h48OJdZRGaQ7NqLX8zxT5hzFfiqHh+/q8+9u7SJADxqftCCZMT1e/H3tFBcraFG1
X2pWNTw90dZ2lK4ZWeSdoWPUHX9l4CwZP9jsvrI6Kltj4iYveNPnZY9joS7KVbRh/d7Suj8gn097
NO1N6UVtwbe3Q38JB7nFeeJR9XJXbLBE/Mn4WkgYbI40BBmn7NsrJ7R+9R2lAnhlkxBwYJKKlO5M
nV9A0uaDGkXDoUdfUGwsOGlGzNAKAZ3PU7IaZNDMF1iPgPY0miLhnYOSopKcDAN2IBauxkj1Ifam
eKQE4h4K44rRLT/utXt1OIYzaS/rfg/FitcxuBarcKOksS2jVvzin3mPtAoqCM9nRGXOCwkqJTAU
XJJw/Xmx3d9IOIUEndZ806l2mJWUl1CalvVtbXGovJ0+1gfEaEPzRUMCC8GiRAR180J/baFrZQtj
zRxztkKvtWs1JpmGrS6CrPbFQyTtJ/40TcoRfNOcDG87IW7w2Y1pGAI4EbKF+GF1iykp8asyiG5I
DJpcGW0dsX42BuhhM3srdBskDoyYE8t5tf+0W5WDOMdpmtygM0CGdBkghhZ1EYZ9nkqcw1GIT2so
FBXcDFelVRSKRXMpOUaALv0OPlaXWz50t9qb4/ZDCCzrEDl7XnSa5OhMNHTEeQpqVvY20tdVEBOC
c620crqr++vWqYkk3N6A5Ph3+/soo+xvtFi09TkA7ZzTkP6UY9KpCbMiA75/rm87XWoQlxlYoONW
ovdZv1JHQL0AEUl3UGcwy1XcP921jsi0vVrb+k/RddQfnVUyR4pcssDSJ2MVcrNJ5lkmOdopgsk1
3vbHQomoWIUcWsaw7OWgAYECdWr57xBFdlUoOJU4m7HKfsNFYthy8G0rrhtfdhvYh+kVZ5Easrec
grQmeEGnV9ueGLwtKHDkgyh8DtluBdwLfT+dTbhouM6eSppAU+XoERJgQVyYJumC9mjfUzZ8ZRoD
qeSwNnu5nva+zzc03w4lOIuzCzqqbuwGIfpBG0/3x6+rzaY87e9ZEKbkQ4ff/32XcUSVBW/ovynm
npZABehXVBvjf9KMsrPGl5W7AyNlJX30VzKw2oCQ+xD3rEOhTZTzgjr2ijnj1fXrveKE6rTKrwbV
JnthSTbkUW9m1IwzFLc+pVAuBrniLlE6ROB3fZojbojnMe5CzdQV3WkCoH/USApr7yqoX1Qmj01c
5Tj7AgVuDiqd5aF3CP0bNNQ/YRPhUWGC2EOXvsh9ex8jwpwg6Ii2VEQWhIO0dhf+aH3+2leGIrXT
fy5q5/leXYemRBXTCZ3vKIsJyCns3kdIzbHRTX6oB8BN1rbxISRUpWEUXsNI8PZdSo4jnZcXXF3S
pljgJF4HXeRg95yVpljieHsH94Wvp0ecpQBOV4NO/HsJ5tZo+5iv+ltK4FHp3+MEvanLZ9M+VOCe
z0RpCP20SkhlW/2Zh5wbQAaJ4vUr8KeAT+wcuz/Uw5xfokHQKStzQA78EdRUtUSE8+wngYyOEOjO
HV/fCWH9m2U5SqxCPAfBJ27vEKeLEwkQYgM0nX7IPuAN1OluhvPjx3C8BosLcvDzffC2xw0ar83i
wdDTmrf+xvKSA/6iE471uqt/YVyvDFeBnwEUNd/L4CCa9K5Eh34bdNwkWn87M1cMvu1BXdMxbs4S
IrFdMItUk5Sw5Is3cM0/8x631SvFTVie5+c559A43vUgIGzhHeR3Squi1Qp0pjFMEINfWKurGOpD
q9ZSIbh3VV+evE0gzFifGoaB9pCRZIW75rQX21i4nIk6/xqOt84GqFJaTdfsjsS7ZsRe0bv3KL0m
i9MWydNFWpkNqHYd0teYqLG7egjYwfp6oiVyGtQISFJOC/DbnktqDSME/toh9JzJxHCNAMCksk+C
w7xpCu9vVyIjZXtxxvWO+0ehHTXJ0GiKIV+6qdltkJ+UrElbpWk11BgSanc0XdJjkjaHKmO96cGR
3TqkafXiTW/ZxMYYMBIu79L/gRdU11Gctk/nUZbwbX3RphwW/Hs5oo/RUqDpn+OqYzBXfP6XK0pz
TVo96+k8n3MOwgYjkrDTWW0MPlr6+IiVq5RLt81Hv0nhbeIiqDccgbpi+HSTetgbCGayCS7Tt/TZ
AMiIC/ZsKmzGrFEAICCmVz+RfDjfWR3ZKqi8Ok6OKBoR319c2IqMb+wEybvLNl/WVNLyzfUAoVCP
bsbn6ggcuLkBGhVXsKm7tEMQzyu/ZjAxXoirjOBtDaLeo/Lg+1E3SuEMis20BIOZZUZIqtu2qqRx
9KBw4gw9qgdEX2l5l/Z1xTHJhrGp2tBWirxkEY+gTjvig1CAs9zznYISrqJMTsPDttsXl9TtDHXO
mBHudpeYLLJxZ3bhdlUs1ECyHAqNYfkWpHknoUGVVyaF6gcrqdeJcEXZZZHPSLYC9V5a4uRMwPLf
H2P6MlFmVzyZWBz69Aby3PUiyHbyUlDRJ5cIzn3nfkZxoNw2lLtnlA2p79ze6k4Qvt6V4SkBm45P
1hibYGIvTgeQhVtOGsvwcqhwh583qWfHCU/k7um2WjPCYM0mBtzcPKeOp4m0cyecccXK1//TLen7
2mrOwLwEW/WjdHpfCbeJdlVIM0O5khBPK7aLOP6G/v8Z8Jvxt5RH1LVZpCywb8KwaFk2XbV0z8gB
qEsfaDIROZnZmbnfJdjOs1cjEnOcQkGYt7i2bSxfAG7aG0r3CbGGUfvwjqmQ/EoDfIYMielkMFeW
tHN9NqWEoCYAmWXybhD52Umjao2SkktGgguEjOWffeyKPe50wBWKw3eVebAKGL7oNpyFo24UiAN9
WA2AvTi4UOc9QXzJgIqPkonfa26+/vgfhyeOp35B/uvFpSUuf7t5CKFrtyh6nMZ4VZLZF/EBQlC/
R9dmu4hmRth0nT5eXtOYomf6tFAUyYDDaVzOPJ4ik2BiWPSGt2AMQQw7UT2ZkI7exlKOJ3rgj52h
pdldpEZ7i5srve8oZR8zHBE4bB5ngpm52YDh5/AKg6OC63p2haVDSgyhcZktln55Np5XMrMzxJoS
LxqvMDBz6IH9k2IU0HS1QFk70ddn7LeAAGGlFFs8+rT6A5cKv8PHKdZu8TTEp9lvFK0LRQf4B47P
IQsFYoB0iN4qQ96VW98XUMxEGnZLf+svQIlQRU4NKknAjr4wFvYBqXBCo5xMjVmYe4lCCnjMFeaf
ghqnfG2tM9NUoSCcRMY+kVaIAV8Ey+Nn1NYRKd8YnjHTFyK4gtHU2safZnGbcjsk3cnzGUmAicYx
05bSmAy3nTmOSsBxwDVmGrTaoAQkv6L4qZaXNmoiQvuqYZMfYMp5ClqPJD3Sw4HxaENA3BtaEIo3
87hdcRRYltTl1G/vHWk3YJ/6kD4G/GHyzSTeY+pSJYbzXDcgxkDBV5rXSvusgGvenVSE3qQHTght
ZPXQL/sMkoiGaUffM4Rnm07aNjz/tA97hc5e5XDBk9KYR6mrgPZGBwW6jSpS5nwdLtQnoekjv9E6
aPNKrTAMFTMrESiQLMH+WQwEEHMlZ5N6BKjtJax2jH4gZapTU5NaVDmde22j90wHLkY6emCbZuqo
lGZDh5XGmQxSU9vjAtCQwICDSIYIXm/yVneFARc1BLivS+nmv1UfkAZ77Yb2B2Fa0nuP8Ihq+/T1
09PxYs3irMxSYtMO/osnc4qTkuwLSDz6FhOmhHqLmZAUDvxboKGHce4qKOLWrCSjs1aZrUIDsBh+
1f6wY5DP4vlyIt/ubyVYj2w3PIk3tNbMGSd1nWEK4CcxEcXmWpRnsg7CCDpjWCXcnuScJJGKBAWu
sMSV1LaSnFx9hhzJdQs53Ogk1IAZ86SxwlhmMpYhEyisVC2bk/XtVvfG8ot52URf3ncEp8H//+jJ
+E2W3jsxOE+STuJyS39Ewr+gz6Uq5NOvdQ8ZafPj5dQqxiH9G0MFNj97Hzxd0DpjYuuqnJMUFGn0
tgmdsNAgTpuVTFOAZvg/p+SY4NaAw27+1LSJYvaLhlzJdbxdwZcXGr+KVFgJYdmgFpXFgTq9yHUL
nT1RNcgnmbvDMh/U+acGVzKW99o19wQIOP4BkQm1cPC8BCxK9cCqcOv1nQMX3rV3QUPiMLk89tdG
t4mZGIDW5lEqx/iyqywypFrQVJ62XmfTHk5cTjcZp7cXQ9SvEKJIO4hk/r8LdNP2AnPuwiuxLA8B
aVwDZGxNNb4oJYIB45rxGjSfPmv3CciVIeII0kw43EVar6JDR2n6flhpI0k34HsZN3HUfjwlXQ7K
cJe1kyHTV0GbpwXTWISeKKjMgf5OHOneO/3bJbW0mjUnmIGP+PuzWFS+29C+ZW0wejO9THRgdqi8
kt4AmDXInvYKtXS4eokRnOE9X4lsAa1XORI/CDfVmpto5Y1zEXGZqc8MxSy1Re/kTTDQZ17t/YoF
C3mLipJvpJdvStu/gcRh3Ku4CDfor3xhaCLo2obxH4bw/hSJIg2E3Sdz7LD2kQPW95Z3MHDDbXlv
Kj+C1ZN8AjNZo2y/L2UF/vljdFMra3dvLBUMUhbRRwmVxvYSoDn/bkOVrlU3EmdyPtHcuEPLCe0D
tsSpDZHY5ofAj9MnJxGqcgzW1odLk2Nf50XVecUDM61OSAGPD4RF30/325EtTKyYdnLLLWCwrYd1
ONf+iXu5YtIsbbs/WwwN7iJx/6CgE3v27zlWGb6NqmwIlqdTQEKBFofd1kvTp5layKW0vqOIfhyY
aH8vURViE6yrEb234vH1a/KhR7bXOXypHU0rSzQ5cTPWPL1wiMzi7eYHLWXFaSTr6XnPx99Mc6/C
3lJKcwnfLpRCaXZX/BJU0KSTz960XT4NXkWtffAzv5Yj5ko/B0Ae1AipRh88WiTwtuY8qtQlYK9p
rjycUtr9VUvk9SY2KwfGL4k7S+P6wRBqbIx1uUNvndQK/L5VOc35evKnN0wtOX5WPx6HKhxRIaZ4
WQLQgenUcr3S3NXNGLW55zWPZkVg7WlP7YdjI8mhr+dpg0mqAcaRXpGaRziIEHb8MiS240sM9jP+
VHQa9THB6b9RJojKgnIG1hj8aD/ktzN8gEYN9flSPJeDXFYTvatQgDC09IyQECTIh7NWGWUMqyjX
iJHmDUx+uOYqmEuRcthZmK8dBMI4BeKSfNJRBh0bioD0q3AAIuIhyqr0mJwLnh5l+I+3AMu7SDrD
xQMwAULF+siWYQdYm7u7VcyNReFiV7nCp6dn171WqvGfPuUgFONsI4vV7iJPb2dsetLqnQHgbjF3
pYd8Bed+UMUDvBPE03tFjSwYv62ZURzGHldwTb0gmtIFbWWsVCJ7J/ocwP6muamZZQgAdEJaHnG8
jfSYA6KtUQhcnmayuRXlbsSNA72Og741OgcgHYEO5KN+1a6IwiJT6HD8dKZN9GZF8KjaFeAHFcEx
TRmYURGklFE4q/4bSQHxBG6/sErvHnxrsfMbVY+kbTmJ2zrQdunKjLqjtbigE2VSSQd0Di7QRgvK
wv5zabHrNg26itYw9ELJrbwdmudCpxdcufr57yO/oEMc6pPtpllSCGBr8iXjSmh9LTY1l3Km3Kyz
K47B2/BfKXTbZ4OxzR4CW4Of3Fu3rcXSVPb/YriaJ2Hm0vBmuIYSZ/7ykhe3hS2BoMkCxQx1XjUe
WPtltbBNTms4ax6xZQjBoEgrF42NM8vE8kPPPLZD2MPayEd199LlXEM72fBH+QXxqcCvbcTfgjOQ
PyXf2s6E2RmvzzI2wnjFS64M+ssKa7Ql3VzF2EXDd6hKgMahbALmMWNe/BQnukvP4of5z8WU6cu/
1c33IRpa1kJPqScvdkztboZPRIZ5splgg4LS464XXFuDWKKJCiCuRaOMGDsrxZWr8b3rzvJmfvPu
N/FUlkts3FAYPa1QvDDvGEswUPN/fK9D8fadYwcaXeUEUVWzhoU0VaHCj3u8oRGO0BvNq4b4b8GW
nWT9x2njBNEDSUIR/lTffIS4+ZzMeQ0iHB9hz3nFgqdQ1bEKRA+ZBEIloL9o1KcSAMDuuF1IsnyG
GRl087OB1YNg9wMMhmyXJatz73zOaG84z16VrbPbAGuUQFxXpIJnHWZBy6HfNr00WalFoTakw8Ww
HrfTo+7BIHTUdy/QNalLzlVr58ffsrao0qnMkvrrTgLWCqxYGNrLmFatySiPjkX2knVCBstZC6vt
bMUVS8TmqKvOzvpkkYGQpdkg8QR3dU0/UL4u/c8KvtbLKkI1q9zqbzrwXeIjtAIyeIITwLlhhtPr
d2xlFdKOV5810qIozcbZN8TegO8A1/9m2e9ULeSip3l5UHkhORVkRcM9KAiibl2VzCjapuyec9Bn
HhDDtCu92yPt+WDrGwycCWxYG4zNOi9nvC1NzTveMnKYVnXz0lacDQ7knIuGfWmcxoioCEFR122H
qlKhxio+Gpy1WCKYF9C+oId40mKsfoIZ3DePjFDg5V3fOleJJ2PxxXcHxj1SXGkLemUTpzp5QeUb
+IyxfLZpPwwGjX/ZDSfpZB9C9UGN5AlT0LosLklyJQV1S3CT3pAjb/saVkEbtfsU4diFSVSniQIz
UfX4NY9hRy3kvR8nHYZucfPN874OHWRbwe2tkDkwRo4Dgmrd2wQ6t9m7Ih42yv3e8XlRe0rB8nkc
8aKpjx7gqHan3D9jOF5FTnvBdfqoa82wsRiRBZK9XjhHBDdGBB5LYspzf9xEnczCsS9NQT7Xq20M
//H/oQTFg6FqpwrI3mzqvVDJXQ+EHDe1kF8U3SOulhRkhp1pY1rc5ys1KOLmFMQBAbTEvvsz9TNe
WohewEizoWmIvXm7aNrVz5Gq2zE4MUnn5frD8/ZSaaofDRdRAladXHGMO3V+8qjNTodHrfipbRZX
mSvV+36f1wLnkhwkUdouB+lENoQCIISW/bDezkY9xVXTOt05D/ynsQhgzpZmlqcIbXS+mo0puQ46
guzPGM00Z52B4QkILCH/Iuf6iXpsv28e0UUUgSrNRMGaQt+8T6/MjqRXadwDIplNJjMXMkT1CXjH
c5X0yVek5aQbn/P/d+K/wqDV50txpApRtnr1TgYyXMqL5nOfV5kWEWzDCzPN5JK2y/BRJFN3galG
tYLOfP/LcumT108xdmxEpbz9iFHDyUmvsxInJT7gjnldIIP0XR2QzBcDsekZxEecWExjg96hnTTl
raW42eOk6HfnilwP5151lFRqmkVuyVr0iGX9U5FA43GPc342L6GVkDVGlfmadTvfHwCwfJF4YDXs
MLIe6oB7Z3kgHN7HpQ0VRaKnf7vhvc9DkvK46NkQcCg69wra00FSYNuYa7pC37RgWmFEDIDoHbya
gNllncCoxhXKj0e+owpkyHEL8i8mpnSrGV4gGd1u8h7dt1FiX5NPn1ibmtQzUX8Ds3z6fqGtqA9j
2b5Gt4EUghoxNPa9HJPAC6TgIO6oDAPu2nd+sYoh/qoMK/bvYI3006oFxeV8KlZNcIAm6qlx0Y3D
cD736cMLUZdCLMDnOx/yLJ2TQJsXcLGg42K9dPyWsPBitdn141Bz/WHYJm6Yq/BDM76wZpHAJ3iY
U7x2aimW6F9pMEivUC3kwJMUGnlhzAEYqUQNrtItLBLaqt4ZPxGKOdAE6eJnDjScP9hHjMTavd9q
Aln2jmFnV3UrlzMm5RRKllfoBm/upKHCXlpOg73auoh2xKSqwwxNTbsZIdv92L3NBbvbpQjanSM+
APKM4EKO/v4ikFxIf30HvQMSvO4lbRsDvIfPuAPV+NsAkFBdiZy7DURXg5zwCYEEPtazjCHmGaLf
terkFxE+J8pDx6OYDWtWwRr07y/kufzIBqSs+acv4G2rmgryepm5B+AmBevr6Ve3S5SFD8pSxmun
9sLnIZmj7Uq9zcx9gyQjju0Q+xz64w+x3QmhP4Aklb3RCxHavoz8Mv9/HXpJFgyCzv/09XZPljYM
Dx8aZN1rleUnsU7LkuchPGdjwpeSgrxftuQnHnD3W/IQ5vu5waNuRO+taB7Wydytb7mOdR3+Bywp
RNA2C20gJHS6byjeLhzynVpwIoWzGvVrnmFxdSDyQlBCtzgQcfhPksbkITZ8gxsaw/D2G5UV8Kty
WY4IUfVtvLrpPxkhUVq5bmsl+VwvKe3EIuVYGAKek9OIRRPc2emSX0Ban5zJOvObQ0eby8X+wmfu
1fAm69khckBVIvwnzA36pUMUx1fdUcCEq6/C/s/XRo/eQzOqznzOJRngKeL970T2VeUneo+uz4jE
bNVx4YGFtmw3ceHm7o0dc46rmT/iSQfDGwxG3UO7g6l8CliZXmV1gT/G7ZmdRQTLsXGH5Ecyvy1q
xkyJ+cyVcB3MTXwZqLBrBXhp5qEYSSXCvdpVCzqV9y0jBDI/XvnVESS+8HCkhL638SoLFLRlNGEb
hScrietKNZu+yMLdNBwdW1O/+wMDjbCpbJxilm6jHFN63rGaVUvy7LNSXAwVKeNcxKhq7NwZXg1u
6CEQ5q0NFXEliBH6CxxBp8epSPlzalrOcFRHCY7iHyafKxZoan2VweHwj8Q/QAUOM1/JJk2J/OI8
ybaWqQpFLvYcVFC7Dd0ZxhiF8KKxH3jy2WEnxZU3/OnCQvz51ohGb6zpEGsJippq6NWeTjJsjEIo
MGTupzdEhGft0rTXFI2v5jq1wjjuiuj1uSZWPywSFH/+Bs/+duxjLAbDtgOyV1DxSd4obNUgJ5Wm
oRsCea0HOY9A9S9MVq5ip33atR81YuKGYlGvIKXsr5R2NRXVDX2WUsRxJ/bF9u1XdRNzAVnNJ2ad
Np5oF7bJxlH9EGB9HfqyvSvND6gCgQNtHCwmKis+Iuwn20bH4BSv7rRaP/psJvuhqlFMd4jDVKEs
F/3/iUrnG6Q3JlzqIxs4aOjZoRJaghN81GyySVpbyzDTaEYDfRTBIT5miBhxY8U9mC3atIVpbt+u
A5yMOT25YkoNq7MxZ0zGjic5WK3rPsE0jjP0oH/WTi/+xgI8m2o8/NAQQ3BoFkx/zU/58EFbtRga
L63/6nzyDNSrMDkGMdRa67AgMllQMNbZrPsDLYx78AQE7Sixj+Kq541b7vxIS+LhuYxxyXmw6x2Q
YG+Kw4IoxOKceEevNrYbXOS3efar+6nTf0LnfY99ckcX5D32N0ZLxPtP0ytbYViKyGq3bTsqsvLn
DRrqjMAWtTSa231FfImPzgSTqWZ6Ox4SU7bRclwsMswP7oP/vj421nvKE6hue59o+menzgakF+Cu
+3bnozRcCeivL2EHM2bVvugeeAuuktsfs2mM3gEnPdMSGIhbbSajpIyGEgkQoCT6KRJzOCZo8hvn
/jHDWDlI8twtagLQvwQk4sYXuMQVkjzSJ96AQyc3ML0jirPQ6xM5jnJEQx9PAxhz0NnuMHzYD0YK
n7cL+cSJlxyxN6wHgg20BB5Bo1F1lb/WgV31HWmXaRj0qhxA5gR7qPWGO32y1vOiZuhXkjX0Pjlz
OcCRIfUu8HBgcz3LpQGGO6dFQwK1OzT/vRNZ5OOb6N4wVfEYJvxCUwcPzhwSZnHNkbQ2KXAieQGC
hwFh8e/PLkffajrado1QwhVSOkswT9BpgFY1Au9niiHpkgpnfPiX3Zf50o5SfCgNbV3hKicDHqed
mQdD4Azga4nXk9iKAYBHqTpnQqh6VkZjTVBTinsm7b1mGH6AqwsWucfzHnThNYzB+9q+7r+cbMMR
ENjR8m5ebaaI6ovhOnaOF8fMtWKHZqcPyRXWMCxE+MCR+L3o2lbwC1r80oXFSOJj35Y4MKVgEUuY
nfXhkgCM9AhMb03gAAEjBFOseNKbl7/CP9CLbCDPVuZ2ia3QhCqb//LT3QQIeQE90PxUwBGiZEXG
eviklkYLVuMdpALksyW9s4zXqc3VuNazMoGh/Og+IhVQ0yKoIi4J2RadkpeALCV8Ro9iS2ZWewxB
0cMGO4BEi4MxmRzAOY901wNub4AiNeDCQ20O7BWpYZjTltH5kmsVAUw0JzMwpzlmmiAKS+EdZ9NE
x30xR8lMz25kKlNTrWkK2/LyMhmhSNinSw4mKQ8K7K8ObPZfe4i9bgY4zBqekAfIB2kbuudB1iM6
Fj+nkm13KGju3/eAG4EvVcCOdD3fyaTmAv9bsigxMuaSxkDkSWCh0AREsfxHwMi38SDOjzU/X9B/
Pjfpw4ANbI29Gi4Cust5pEZ+zh9ZCrVN00VUa4qyrgMtkt9KdDaGTbpPJbuRXCAX7nJqnawZRq3z
nCa0DT4a7YJ1aEmhDazaoizPEaQhsIJKDuVqHhPJ1pKVGiwicYgqxKJtLe2v1kXnan88SpKuHv2I
oB1RE9kAEv5gKoCqz2qMc+/dPpXjgBYXsQcp+VLHKrj/KZULm0ikn4LY7rVniw3FAqVWvlOnNyhZ
cwM2YYuSndxtMznktKfugKuLC11czXlYyLMlKRga6eUJlkTDrip5AwQ4lGUgbRFHA4W3FLPdfXbV
vFMsO021zCEBV/oV3AN9acHfpWHd1ctFK/ZXmQ7Q3R7KDkCZJbJskJWf3jQ6UYQYsGrzSbi8vd7q
s74LUsPUcUTRw6zKBABPjYd9I+De7HIrzpmZKuLJAwjR1Ppiq1wYxN8NnPW1kpei4+GUb5Nm7yNg
rqT/OOlBGhoElKpsYUVN0YZqMxT5sXck851Ey/WzVTBHq9e3EnErQ7Qxo8J1dY5P/7KzHgSVi7Lw
DS1rPlAqCKyc1YDvwnGSvbQi2B3z0P1HtCGUsHgnt/Rn2IuKXPrCxYNWA7S9Un7bw5z4wHlPVTEX
DmxRnw+riJ6N/gPDBpfUeHmnz8P0YxPrI/wYfAxTdm7s5Tg99WWfF0f+mv3ZNcg5U1wGbwzx3kIt
6BiVGpjI7ZTnTgjR8HEaOhXNgLZ/CTPzu8zTwED/ErpPgkXShydjMSVXD1/vCXpyWXL+kIGahikV
OfABwinC5aWhewB7n+yd7O6T9Z5H0Vu4PTQhmBzGbRUVySEZH//slsNCIB0xeONspQxMUni974dG
KhpcSoLZO4HvzjKHRsdNhoQconOMBSP5bWCwA7aIkUNeZv02QDJ/+/XXKQ8UNGtNr9lDSD4y9gaR
Y0mHXexwYzRjD5+ohgaCx9yKukO4zXBvvBYisVxyte/7dhCVdGK5L3ek0CDreD6omTCUy40kznqg
ogm8mgnI0p6QDJbdbChyXDV6k1s3kqxWu4tc6P/x6hWhcZ4+yKcAgHxT+wQC16vkichy11Fwc3Ut
kz0DoadJ93og641k0QQLJ6Uo6sLIJIudvamrbH2s546B6JTtEG+tzLb6K79HktBnnKNEInJ3ii+T
fex1ONu6exKrxn1jABSeZK0qUKd1ja6izq30fUADVZ7b7Nk3huol8w/f7dBrF5HeP652+TZjA/F6
K4ES/zN7gxREc6hNJUW7b9Uv0uaUghQx1ttHWyH+S8QsKSgt/va0OYfkrkpM8s9hmpwyGBG4XK2E
8FVs/dDg0zt0E32TEsmILDQ5YfHL7WaH8JSpdatdVEk78MELt8b9UbLUMooBO1Fy6IJoV8iNL1Vk
dDjttvPgKAHZkhhmw38tGAxZL2EjoiUoL0+uWLsMS7VER/aH80lYUiQf97dWHBQbssMWXXlRl66N
6Wq7FXYw6r/WK+mu+OwdD/vlbnSN/amtbgwkzi7dag3QPvUMag4ud9+8SyaDGsYpeTtoFIE7OvEJ
Hc35tLDCahcjnoF9l9oCMs3EhyOxsqPGBz81ugF3maeCaXxI0LemDGLMN9Noo7VMLOix5TWFwEaF
27jTi/bACQuqJkMhbt5WDS/a3pzII49/HGZlBxSGXYl/yuWDtMMcMnox6yzlFRbiCE64DnZgKnbs
z7AYNpYMsaPfkwxZ+vGcVLzvZYa6iKD1WVdMce5x2IpHvWnB5FJFS0UrbpRz/0jstKax5lM+VtYB
7srTFBj9qLICvjIABYtl3M4qTGPK3uR3XbXxSlW3Whp+4z+8BbvP7Br36tNlLm4Pq/SLu7r10+8X
0BRPaW4jh6/KoGr3Xcq6ggywqhMbKwmhSVnEpNPPFQ9yphowwAaQ08KQl6WK8irqJfsFp/9g7ojj
zbaNjoQNMOf2xxPmescpJPqdVwU92uhvJXNGidYb55qtBhwfCZUy4h8tHdnBw9JGug8iaUayocyQ
dz69qIuewXR9IMWGexNZh+/F6g7MtKkiMNAv06mXY8dCfaOQXfX8dpYkGw9++o504dsvC67aQE8N
BaUSvPUfJSIfdLUgoLSpt1w0UJ8o+aAQYqj1SiBmd03mmSbi7xb55OF2psf6DCdXHQN/YI31Otap
QiaxYK2p0IyggPz3fRE6L1y5cqBShBTmhnnN9/okyN8Mcy7Oh+MjdsSS+6ZF0o17eQlpAv+jbN6/
469EFz6f5cG+CS0EfwSOlUfVJ3+IKj0ahP6WIyihl8ydw24TDCxJdosXubQ/tLUrlbrntPtX9xKE
GoCcBdCqOrmotVrhjpqZfD1KVgNgbNXXXR0sXB2H3alSb2BfQqKpPLK3YcIolJIPb068m/FPx2N9
vqtNwko97MnnSJxh+Yj85YX/Io57YC1v4neFs8+J6Wx6aCzaUfwdOvtG6uapcKd13iDOxpE3XOAi
1cHFIOtsuE0XdMidozZfyJNuh5ylsTAWmyBbvhhYkB14ZFlEXhnDT0x60dT7/xkDDzOK+AbnTKPL
AHqwUULy9xy1nRzyXMtuYnK0zejhzQbjcH6uCvBcT9lfS8Ze4vYfD3FuIfuoUT7vk+VX15P1pz8K
h8/AOsw9e7dZLrLok+3j49Z9UfvznRe1xgv6CKzTPW79w3qrUm0jwrjA0bZihMFMA6E4sjlY0l89
v4fh8dsy/oCAu3EBZJ8hQv0krlS65tisQfrRO/ikSWnoHXD3bCncftkpzN+hCPg3eQEzfCfJtugU
KoNSz1Q8VUmSYTOz4G+MRvR7PbW8PkG5YHNBRT+L77xgRRpXNMNBoKss3kI4cNwX0ug6PRoWTsi5
hJbYpDOK9Caq2u2k+1VF9WVSxyJdFozvVZjuEqwmlNNl4PPgMDVGXQOsIMA5XRaQxzIwjWy2b8G1
LnSYGuIKvDJdAVcqYqd1gytWlYiWeSdTB834jhWA7ox5eTrhHH6WyZstNV3GK7R7iLlap0jJBfpY
nauaz5kRN1FUBbd5PZSMy+T1MvCV4yuYNyBcYWQKVf7ksVddBOHEWy2njwg4iGKEH79WPhfLszTq
kNZJYETago3rbY32Lr59duLiT1hUB3lsc/1AUuG9DquzqBk9KLvmgIYAYgrg2pyyClE6k3mGnW12
LP/aU8ADMWzdzLFISqU6zOSYd675KjUdnQLu+OhahW1tk4ETdZ4Blpg/fSUyhxLyovgYZrb5wQtb
rA5tHKu0lxDxv9GrVWPkduJMALBdLLwGSLUNJG4z854MZU+RIpEzYqNfUJOrALj6aMj7ftyJyAz2
+nY3MsesgotRDsQWupTmDc6+X0pPFpVOhO9SfVIb1ZucKEqTRy7DRYLERQ1nnEnuRqmcizKZxKMH
fGykoVRBEMjxfw/c0Ie6sClZgPrSg1WfNhZlhCHgwUwIsqIBkx/yaxysNT2AoVo+NpNctYerprxv
XWodT8vz4vVib6UbSPrXEPXquiSVFuurxn2FHtLt7S6ws4zDoLCJs5xH0uEG43JTZ5y8Us44k7Sk
VOwTQgqwYSS2OtGZD0PpnMUgmAGwtQjbHc4T1cARMiR9oHyM38QftGlK/XU4gUSGumo7RUEZR6Up
7ks2oC962rbiLrOR2MiF3pFs1X8+ECuvG07O74MMINLmkrbJh9hS/IzgPmqHT7VX2hilJmE1Src3
IkipcVyl2N6mKakgKKLIvbANI47/Ea3y1fL0wQ5MHih7MCQKJs0WQgRAqUCqn27UIIj3HHkfNoUi
0vFKMcdFmQ1RzqqKAnN6gP40XFMu+caQai63bInZ8GlCIPiPvApcVSWFB4GCxe3X2akOiuBCqlh6
ZG7P5pRn40V4PngZ6TOpoifPK5B5Qa9gGpvphKP1agEn0+dHdBdJL2ofq02tz/bTtuDXpCFYy6Mx
E5d2Ul27cZeOBUuOScMraxLRgR/nBwrK0rnPLJt8EkfBM+Lwcvsbrcy+3oHy8Wl7Y5xmJdqy6/Xc
9aDSBrdx+4mklvdnblIexeDB9Jq6XVx4aaNuwNnsDfPWVNsHoKj8LFk23QpOrQB+d9ThdxYHGivO
q4Rvlj7rKR0tYanmwbUzxjDTgR7FktFjQMswJqD/qePvrMcGFRGe1LPIQ8LMuQNyGh3GAmTfbC3O
jAnn7WqpYkzPyPIYmattLqF82CyDVRcY/+db/LCd9rpyOFcjjWOXQY87YG+9JLES6h4uwYYHX/dq
rBB6QWQlxSBe93L59TtQLa0f8AKg66M7vQbRtjDn5NsUG+WfGkjXCeqytlbJyCm5wNXcAdbrJOfc
XeLsezfsLOopwW/wffTcbx/+7GmreMPcVmCOk+rqrXauu8VBbJRBK2PKY+9Sa0a+ea9PWdbNKk3Q
D/lOWZzaA1btQiqewMrDVxOSGN0MAIsAlfmxdr/OHTYTTtErvS0wDp0WkN1BwgK6KwXOpOuUtCVy
e46ti0w/73dkVgukYbpJWoj/r02uWmj51CVx3XGHQLNWhmRwNeS/By0U+i1B9ZCTx24f+nGHhuNe
80MNbinU5qHGPnKgQFI9vsPF2c84jWWf6XIxseSI+HXvAldsZjHYQCE9Ut1Jzg8GsmH0IKgh/LA/
PTiQdCKeQThLZiuVZbscuxMOKsZAF5hxMPOMhTiy2IWEhA+L7EJ0TnPBgBgAXwWOL1QeBcyX0j0S
7pTxY88/oI11X1lRBzj0l5ThdIM2FeGO7xMZWPi9wj37UopSbSGz4Sqi13lfW0OYcbcAkfx8Hxca
Vyj/XEU9gaJ6OWosJBqTwyYpoLpl+ofjmvQsUxKx3za++/gA+7CGZS/sYR8m8bMNwI2EWEmzt29F
mnXPTQp7ZqOYSnLmHy+yd36TGuCC3Xyi2tB4KplLZL+ieKdc/rSVT5jzcosqhpOToOKiSbcs5p15
Bk0oKnV9CgNgQMfA8C7xsZYVq4SjBRDWYoqdYnWDmT9CbLa48k9DoGXEjJSC2wAbuX2Mx2I5MBAd
J7OanKVSGeXhjnukNNpVEpKXELsaT4zLfutcwaPUWVKKtIQZLoAqJvg6qbTpd7W27qyjbHQ0shc8
/ZYrH0fev1M76FCPzaQVtRelfZ2owxIE7etWUc2FfRhYd4SmCjU7aag3efv0mVYtfUJqYfRBhozn
tjmYUkseCwzzbcoCyDw5kL1ftKCN7ND+o/q9t1SCfxIzzaxLX+LNUpPdTNQG/ziAGOoSUsVz/0tP
1CMPpVHMM+ECKKM9XZ2YfvgU8SgvmjKGpaPQuXdvmzT4GIzSWqs4UrMRGBqp0XHAiifUk7j0HzUy
M7RgQP9I2et6j1UqFyK9LJswKiN6y3hYmtKo52RlKeiKh/7m+jzZSZSRJolZnnPzYRuBGiseAkjj
BEuPU/v6N3LkFHjehPRvNGqTJggMwkvB5iIQjf1LdniLjaGBc5j9cVrVHy9de/l0TxA4ULOV1zFF
U1pjUNRXouVQmNN4p6Aq/aNKk2CtQPwkPQhjUKFcABk4RpoQ0RgttKvMsBhXxTFv3uxAPt1MgT/x
ADET9pVRmuHpWjoZBvhjgmKZEy9p0DSTGHDQIOOmyCi+yQDVBAZV4dUjWA8Qe/A03TY9vDF350a9
povd9BmOqBMq+4H3KF5urAZd5O9GtHSNkR/6rQF+4OgwqNXxtcoH0yftSVDwvl5RwdgVtejvAdO9
qVDzhv8oqTHXMcdxHca6LMQHRrc3GDRrvwTyH6AFq0qV1GbO+KMsJJoxC4kTKba0vIMNgKwagQd6
+0s2jPPhkjQQ04DtM8ShmCcgwJRpYoWqqPk4Un2J7P2fn0//pzbYL0uhMttrxAZz3HHqkgr/V6fF
/A2uZvwrRm1pGt/6mvwrO7RQOsFlyRO0PKwF3ak/7ReC9llCqeCGDU242FPriS28hQvnP77qvR00
yV+J8RK4f5PEIDWlwS6JFsY3ZHt1uzMd4PGGhNcMVHX4bTxcrXll26jIoontpOEEO0LSqEC7FsNr
pfWDo02etFSyU+vNN4FUlKkkyK5UaDS9PAHslGsd1r7ezTw5OceydYMIazluxO4dq7mvGYtgfpO+
Yew+fvh1frT11agYSLLJ8d6ZOlv8REoHb5iDYYex1czO7MlSUjP4ioIkFg1WiHtywewl8bnOdUHg
l9HTfdEAjDo48KauiifO2zR30OdjrjHn+2Q5cDpnI4Tu2OhrSLzFcUB/tTSSpgd31Kw3wMShwzzE
jG769KromwlTcrM9hetrD9Rpz1qmNyZlmjMZ/vlun/clKM8ReVlkGCn9bCjLpr7MgJyepNwDd+lI
C0fVDevgV2HEXhWUYlqkn0TzNdrChydX0OK4E6EPvxg0m4jywn+QtE4xfiDLBtVmktTTr7GD9/+W
yXAbJnhJjrCvmwGzT8joN3fmY7bKAwk7jZd6ZE6JWTCkHKvSBZCcGCtxL8VoMBpIz1W0t9pnG7dU
w2b3UxZVwGMaNlD1peNywmO1fvPUjUXTqPvQq5QmOIOJ+ORfKVfiiAwMy0c9Pnns/tXEF22FEaZb
/M/JDe1aui5ZgYkzT6C24H29sPGSlbBBTiXsPI4mXvz6Taah7Qc9+ggNxzt5YLmYRifXD2qeBUL8
1J9/7M6/YRISqMPKAt48HMKttEq4EizsIGO0tNIOpJ8WI247QtFngemOyrJdd/6Bnv31lE1E/up3
x+TpM6vJKeQsLWeWqMk920tWdJ6UfCWRj4v0iIBQ+LdoZf/QuD39AFHg6EBT82N03pNY9+bda50m
2wNEf8/pT2h6S5PhORDr0m11Ilh0MxAggQlFW/rzmXTHKDeCWD2t52xUZ5BOYvUlNWa/VzqyY+BG
pHdG11M6DmRIG+IeW/DSrRKQTLXDdigMRsyAxbiyhRGj4Z2gf6hefPpqsbznOQugyo/3ILM1ES7w
QUalW+hWH/6J6pkMQWmM3kUXrGgnwfYi9h0aFXGy+W9T3o1KGO+G9uBYq2CG0v/6LWyH6CYJs/Zh
pwxDPxLgLm6UdxaxfgIP7G2GbSCgY7LeH7KH7tNxHXpkS4MbK4vCxQ9kqyB1NCLYzWBsLLszV4FU
w1SGOwcT1DVNkOPxXKk0AF4G64ZQjx5ExI/l0jwdmwvVxObCULrY63XC+yX83znjveIbH1WDHHD1
Jd8+xYnSLDFvE3+SULSJ+Osnecw9C1Sgqv9VK2sNgCGl9jCNQ34Q4kJivMkk4RmzTpmgAKSbNyvk
LLtlTUW53UGWsfeqw+/S6NH5oY/gvUaY7rl21fE9Lv90pkC4GYd16xFnr4KxQiGePllzpYjDfdTn
CpR/dmeduDAOdRB25Sqr2GxytOH4kQjVUl7PYCDXeYKKlORBgT4kHRQzhlEayDwz7pHi9Pwg+wlP
6Sl+hO74K4g4KGluzP2sW0AktMoldrlZOBs2U6B+KU9l7ngwSUEQeBoBtU6xeru+wo5rGrNiekeC
+KTawSq527U1AF0U0onAA+7Oe0UMxv43+xxE+PAtGaPgcttMiswMIkLgOpg5jC1K/pQn6r5+ZiYi
i4+e/aw7oYeM0zInNyUR/mdRyluzHXOgrycdkBAeO+rDNafT5f+i5vgf0hTbqbSgAypWCs/626KP
68H0mO/TF0pOkeFTHZTtx1lY1u6YAjAaqNvXzrHdZ7ooNlv5z7JPJ0f48HMa8U/fNhNRRTl8C4Oh
K6fAnC2Zettf6Gmrt4VaBEK2nol8R1nAMxalYjEiuUOQgxLwnQYQeU5ytPYW+tlvdn5I5bfgp2Yg
r4XZma9ONrFu8Z4Ekp3gTPvm9ci4n/X3DV0KMzSrTB0YUmVsIdT8d0u4OfsMRWO9ICluNKFKS6A5
YRtu1s6eNWqG5SxGYTW30+ucWNK4u6m6fa6kPiLYnGHdiNN0F4EPt3o94ajJUT9m14VsF+0nlVp/
1aa+1405Kk0+wBSbMsPgFmc3Kq2Nq//u9irfd/NW6yqGSZjDCukM/U0g/FG8XYHYa2bfi3J9EaVF
Uk9zCcBwwFPsSB0IluxVbiO3hAwlDvQ6Qe6yaBDQfxOVBJkjXy7NBtOfvTIfwOVJ5wJxfYErWxJ3
MDMqZZXhqIlPPOlDBB8Wdf82G5LXFnndnPE5wfII+6DhK/KYFiuCaOTJqykd1NPXHqx1CaCoaORM
jvopjX3w0ubpgEugrUK3IcTEVtvbexWoqbrqhbpMVD/2Q79b+JNSK/d+7vnjShmqzPtn1lloIiDB
/mDpFhmd6hiD1LUVv87OxebF2V1O5aJT8BHn/B36Djs3XV0Hjz5znT1BlqBXwoumIV8QNRHEktiY
Sa1AQ3IIXJDalxYZzYJeq7Ky1RFdbae5M3ZGQ+6dm/CgAT4aatbMNWZ3SI/c3jPxsWA0T0iawrRo
bWs6OLt92bvLv+IoeXDXiMIGe+EDhsuZaAM+YPTD1eDBVRom4qS3er85WWP2XyQ9z8e9Ckik1Loi
UyNic5LjxdeurH5KIqCa+LQxIEeOZ7rPfYC7DVSavwOLBHhaNgDIB997C0d/OBm5obRSVqHVvd2b
AMiQWx1I/oa6Qjxw8ofxwPq0J5gEpbavbsy+gJqBtAb1DIhsKvjexcdrhbozxcTAFOPts3ryrfwe
v4L0Tcy4xFY8rbu+Z06aRageUJruzwg7RMcNNjyEgA2wdTG6k5GWEgXlEuzivZWcMDbcV3KOjkoh
Q/dd9Eh09xZ6dSdsa+G2MN63Ocj/tI+YhCQOz7EuO89CcQbm2RvVsyGTUVeN9+obnQZ62BZ2nHBN
7MHF/FbHbovXffU77LwFEbENwxzZnog+PdBzST2TDoLmadBuArjY/28uhbyg6f6GDAYrfRcrs0uM
5522WIDBysqGrjAcuRjK9ivJyhpYJcJSdYpgvIeTWm5l/rdK3HVGWwyp5Awq0E/HUUEpStLv56Pm
LtoajNdMAQP0xMHWImubkH6jKyG9ftE81Q2rrEHvsTsDLjPyBK7xk9lFlPtda2weNBet4a1tW9vU
SLGkANKxE8H7g5cEfsZzYdhpe9JbJylnfkJLqMnPrlnIm5qI+a0VZ57cRyvbVqjhWeMrHIvJ2Oi+
QgVfujJiVbPWXl+TxF4D2uxMM3U95xVAdUt6qTpK7WDGasM4GLadbYMPNLezOjBPcofWDsS5I0aS
cbHrZ6ZXWaSLC2SXVihVRlJWHhC+UJL90AbpJ4r2SpBR8aWrp+3t91ikMAqWVvmvFQmsvKVVIo4x
mjqQf/SzfCHPZ2SJBcXhh5dop5eD4PC6WO37trq+GweAnt4K7BQhOxwT97gYAAAp/ZG79yc8luFb
Mj/FmCAx8ACu+wA+BySI4Tq0SaOZe9ginyI9eYSNPfTSjtZWf0DXxRM3aPhqqXfNx19YAx/QOVlv
hlfeSJzx9UVPiuv5uAvfThF5Dt8hI4TzWZUh+P6BM6hhaBJdAB8lNAEtS9Ftyix0wBlFxFcFU7dt
Vz3rbbl4BNZ65qzO8EiIqGRwsaUvFNR5kRT4p5QmePMK8pD0aixJVDFT9HDdXyiw3rO3JyxzDQeD
/dosuS86suBrF0gpfXgYbKXHqJJPJYZsPYelZBVLG4oNmnIxmdEOOsCVyVYomAvUnqy737Hv51VT
e73xQqfBIhFZnY4IQtPLUMoUoFAx6lF+leKFqb74DNPLx4w2ysXNuUrKza8X/0JEUM+YqxnV3lf9
uZqm/FhUJxaiq4zhAR6LUu+Nqw7VJ1n78pst0nHd/l6ESQCfGRrtM8drP+Xr7nF4qEYc2xKunh/G
TDdRJHTKbmnYquV4ZZJNZaxL33AcGugvCG7YEE0r8wPOSDPL7bdltEgtnePETqm+bdPVwoA+EKTq
vg2rCQUiOwosXFM4Ls2Xtetncbp5NcNxAJAvExXozYUsXCB0BrkMAe7XavrFEKkEfaw+lApmxAJL
KGNK2+Nzq2Pk5Hkc6Tg9Z+x1R9iXmcDt/i2r5h3QU0lfPdq+0qEkBRQFZbEpLZw8A8GUT9d5vIOD
rM/rVucG13Kw8+/gP9YbyjVCtZdWrWoq+5/n+igK2RI7SsqsSztsBfoyfLw60uTDvwivHtaDatmi
ZnHukrgqIvvhLqphIILGMfbaY3CGCJqHQqmXVLc0sB4/Y+UfFZ8em+mGTqLwz4naQ5bMtr6l2juF
FG/pMyXX1xoZta3lPqTYedEzeYoDcDqVO7UcJX7lQavn3H0PgkZH0cIMGqOLtVwcHs0/PE0WZ8fM
xXoKLPQkoaHYo5J2hOlbhhgGpBUqtZw8A2SmHUspEzr19g8BKdSjDXB4m6BFRB8dwzY4pbEpXPib
7y9heibI5nRKpPkPQnZV815HTlCoD5Tydgwl5beNJho/zjZfI7ke2eQlxbljBE9bH3QoqKBy33WR
kFb0VmFbHr5mJ7p/+sravl+yoO8quQQRDmUrBW9PuGUOSv9KnX1boC0qpDbhU89bWBHb53gO1VD1
nWZA5Xii+bIhNxwJOAmju+1molPsncd9yOqxvkAXsY0efIXBHPG9HyE627+pPKvRDgbH2mLvQHR3
ynmp1/0O8NT4n88lZ3iC8P5IcP9vBhdgPl953LzIXq+cSjvQ4Zni5PbSjT2AyDi3LPujE8hUbNNf
wfYi+Q6V5Ox+XuCmC1ko1MrECy7sqA2i8HWPLTRnOf+jRV3JuDp7opAhcwqtOdIpU5s0adDd84q9
XJzE8DQikW5UbkU3DYeRAKCNSmK2/Z/MInIiUv/6aeijYT8Q1qx/ECibm7iJ0MlQ+dhjG/d9wzVx
iYX1zY0rXUtjzbKUPyMNEhqHz5Kf5nalPK7S8vOw45aZEwZWUn+FxsgJQEkSNymmMbZ7THRQBgkn
/XqgxJg8z2T3xcICH/ILVfcAMEP6uD7hY7KH7kg7pJYKvnF0IWaRMROcR9PihoUyA++BLrw/4Ana
GUsmR+va2pP4wtDJ8BvdzV/kDpZp+hSPvv7njGPzqqkJiCr2piGssWlHVfaFgm0rSC8kHaQhYnHU
p1XYG4yd7vQ4HfwEpKuG1Mk0VA08lCYQQ/qucyARblPAf3/HTBx6G1QJCxUtWWyZZIP/eW4gnzKN
70N+hEQd+AXnOem/Hry56beYp7an6/kHdLzZyfONRbMFHssOpW3HI5YguUxRocTgX7Zo9KG822mt
aiByuV200mY0jMAB4X0xahS4dtN2VTCmEv+ieMBk1EORHFBryoM9pDPX8Kn72Mw8oEx/u+dYHg/0
JWXJNAyIzZ1gj/oJNig4M5M2cUmJQToE6xY8PhYymPGzsBqsaimji5oXigEy/QG34Rf3DtA4Lph9
PVeui/8wh+AMRxps0Lo7mshYi/YilzWJdObjUmiqiZVwJhx8DwmNUXmGzyB75mHYMx3so2aiCIlE
oHbytmyOTLkA4OjIwMwE94pfnRvQAlDD1ASqlH/CDxmTblmCAr6y2m7cwnqiKXf7t3ciem9FLNp9
n19WqOD5jlOSQQhJ1WqLxovZKlNBeX2hsS5FA7T2qmXaBwrquBl+/Fmfw1HeS0jFHR/9gfl6fUvb
3eOb36uBjmTjpHdYHCD/O43Qh/HJVFbANrzzQa9HfG6Ws/0QZgGVptGr8jGd8LK6JuVsXkEeRD62
Bgy9qYgf3NqDvKf8ZwKuVfIEKgDMuzJ1jYl5lFkgdrfBBSzoyc7BhTJJV0RVSaWNgH7l6BCKiMhl
EoJcq+C5DaVLKt5eZ7/wSDXjiwiCoS8cJjYB9OC3J+tvdwhL+DC3QnB7ktBwfyjWJGWSWqEdWWyM
UYY4XvvtrgRZXfQyIQXDyRttZLwM37L+7GkW+H3y6l4cUCTqn5yjhn5XnQNQJOkQ/2USE/IwOY6C
6bZRwxtnwG/6xFlwZS2iRR734RBRDhe2lHc9jNaNgSl7NgBhS3sbZ8m7q3k9Z59+BYq/V7XkFzIH
dGiPmsnOLC5PlMPEDwwVbM0SYLUcYEjx0Kfg1W9p8SsS2XHIXhywnv9RlGepwfK+hNT8ade1uMhY
zMWWrP9Ultdzg6gCZ81NNu7VZWvLtH0wcCKw1mTGVHcd2DmC0MZ9uajkwz80bs43kItWu9UFLRxs
ygAE9IJMwAKhQA6cZvg+emJRdplgg/xJtRFI51/XIMaSvnEvcXQ2bavbd+kDLCWMzRIxhgpGqx4v
joEwzCqd7xqotE42qge3mMWeOqn6k3hKBjlSubZghouqn+vV62aphvDfUS3In7Iv8YDG0WqvVkhK
+XMaTx7DUWkNVFdXY9w0EkiOAWLkOAgcO7Jpwygh+8uP/FOyWW06dsP6Qm6cvjx0jlUZ3aDe//vT
NyuA8W6rrerCtZECRvkAtmapG2hw2o6DX2pKokFmX4uK5F35MYsLd0ng3A2EBlxbx2KHuS5xZqRO
eQ/GeAevfMGKrkT9TCBrzIWGM4oZkb7yoajMrZ3YDb0ilEKZH/BPZh/26vEBTXcuQXUJ9c2uO2op
Vn+vZT+J+AeZJYXsw2IgbwMLkwBt/Pp156U0dbW8XtzAkglCluqBRdnuTndDj8QY88cQucr9ip7o
xU9n/Tf/ItC5Qv73Nl//ZbJ5VDNIzPHcNBvVOGsYdtHBnqeSmNYJC2lAKFWeX6QrNEpvQor4I6IO
g0XeohxbKOF8q5yhEK9iUvxxTtejg3wml1m8bsfstjBHDIlB/zp59WK0rspwjrflE6SQZF2rJAta
xt00fSpagoKTe4vDen4TtLI1incb/+AyvJidqyOQIfNcK4seJSILKIKYRAyBXJ8wSPzSa+NykRSc
rzLh5Oj1sFjKCnCvEzBUYP5ci0z0zEqQWPnG8oGwCIKBlAWk613ubFIGozlXGov0fQTdc7ojVn2e
2y9aiCQlcQCiXDzopjvNU85l0/yjqp2PZHEUh9rjHTlrIFSQ6qvgh5G7NXC+sdA+MqOovCQB6aus
qFO110v4QDftgpS5l60pqPY6bKE7TXH9RSRXLTFfTBZlWeUpEh6lpGCeu43GmOy2CrOfgIX7uu5m
4rBcNThM+MPLPeQvgjZHDQKalzVZOHUbMqzr0NddnDml84sYXMH5SouUB5GQIwPN2wf8Bsr4tMpH
/3ixM8hccp74azOtOGlo/5l1oxpygS2JLFanCqg0i1SLm4SbdL9Z0wSNf44PHtkBZUzpvxgtXyU0
uxYNfEhZDOMzWtZxxYg7ai581wdpCDTKY3MxSTDEeYD9MR9SS25pczQNsrAIVunDOMpwTeKyku9B
TxOJU6cVYonzkZD7lDYjstee9qmd8pctYvqT7C9Aiim9oppYBCrscxYuUgPyZKRw44a9nbJt77YX
5WBLI4xAASQD5I8yTDCnHLgV6V5py6rEjIhgSRUJjHqBSIlgIBEJvRRelwVmbqNmOZ4T4LUb5ado
0UyGirpeQjLL8SXK5kxVJ9FHa6VeXuTHdl5l5V9YDjEbfGh9vCYXvqzFzTItfe5byfGPaB8VoKnv
RJCwD6UbiItCoLhAfyu6+TgX68IGi29YJ7Q5/Hnum1LrQqAptFGEJMJkB07iUyf8AS7MjuRQ+ya0
muitvKAxRm7TSUkjR8MGTV9iJfauSIwm6jixGHdujFlJG7r/45nEgOQuPPxOdGR/Y2ihNhpYZTzW
5rnyIRcZHnXABzCuEDknoOPdzMkHrh3CK5J9Gu48CGrEq9jQUgyHK5i3Zsz4xhgrTLICoZdMNGTQ
0EFctQ1y7jTCD4fOdZeONIHICWX3tU0WsMHGRBl02sUvyBHpy001TB6s9OORtZmkR0wE5jcH8n42
I+9ab4RdWcbqRdTsopiXzLUvDtS89OAXsoftqREOyEB7F//rF9lhk7d/UynCbd0VNMqwyMvBBPUo
qbJQi929olIwb1MqIz/xNAbutNiEjxLcc5mPFvv0sGwMvu7QrPYUeDY9ugObhrDEscx2uK8IRA0F
pt+7G/N52aUV/qkKrsvxft/Pm3nmYFKCnROS/jkpudgkXgAliWNxr+xW6penQ+Y2qatvfH3jVTze
6yjUFA0Me73V/VFzfZ8iYax4craw7O74mhVN15TIqMJ7lQZ0CuRkUKrRNQRXK1oeULJlAy8D9rH2
bTpfl6kjBEOav9iGtAlCk8oEaKktSoLybD+N241XelFBxVgpIQAPiAkuXmyuEPxqUKMWuvtbFDdY
2jNy2vCqGLvjNWwez2PIMualsmOjF47bihvsWssVKYEs1enN17MxnT+Dmi3DUlAG7Cv/gtmTJsl9
dOje+Eo8kf2zCgGL34RS9DY6wi0MzS1fwkYQWni4WV4dxL3/8+q+TIpOMxOBtM8Gn6Qj1hiOfR/N
4DTbmEDgwIgkQOEeeP0ujQbmTg1feOoh0pxFOF1cLiS2FekgxsAE3a41xm66k5B7clmJ77C+Clii
MmhvCBtV+W2r1FNuwm9LRXqLFJYs36DaOn8vT13gdHoaQvPc2opx5vAaw9Frs/hN8XcGapST6dU4
EdOsHTxXyfsU8JludzkhkgoJauIMAWlYk5/hjjHqQGyjOjrc6sYeyFjOAHCvVqzJIuCmrepJQKTS
1PF7gwI0T4ndBK/Bf7VF7JM1RLpFbfJOND/1VTopNez0ykt5Qf9Q//APn9cLMOBE++Y05H4SlGqP
kTlEao4n0h+843ebbatkcyIPrW05gRAIGQNW1knvPK0MnrFoxAtuvbEW35aDoQc20hiBZuyiVP5j
zldozUVrla33XgZVaOjWGJAtfnBIf+dZjjFKZjelFZTubmULAN5fzl3M/4Z51fOXiGl2/Ny6HIoX
4NaaqAjJQFmfK1tDgBNIX+Ksrk8Cm/fEyLLWSgikZvG/dpR2ZvLBJPZhUrpEY2K3tL9iJdyyDSdt
QqGt9sVPnIpi92CSluUSSMV3TwkVb6mdfrEXUB1RP3hkNTLtQk+youLZlJoJeSTQcy6NPTapqHKV
JQ02pYgh+ERcuIzWFze6VRo0kwJKyIjrLfkzOZsGbidrhyaREaVRP/v66Az3nWjIKR5FZmyRFRXO
9ae+AuwcsP/ACDr5i5NCap7BF0SNBTkZ9SotC1zVwNrRJASY3EUP9SV81yrcZBPMB9MgpbVuK/SM
3zJxOLHOzJKYcblDtNSNeo1CRMH3Hoe/J+LOr9BFZUKZ+iMBZ/GYGPc/kEfN/59V3BhghQ7RpHK7
6ykPnIOpCYfy5L3mjpqpwCV0b2Alc4fknO6uSoulIGouOU8RRO5+DVjgANkyL3LfdQpLkUJ4nxeE
C6OECQjzicVGWYZ21Xsilqos29Ew1EZ/zDvzcMNptg2Djfh1KydVkldFGnZ8dzWukEy0r+fdlawQ
Y1F7KhVIBKggpE+e4WlvijZ5sLwBSsMBQF6C9CeZN2i86o4iuedvgIzQWxzf99zZpqehK4L4IaW/
FnTkMXkhizzHxImKl6GPzN2hMSQrFAMWvy5KJB6V/AK2bXo2AEcTAfRpYarMKTYeZBuIKcEkIM/p
7Mc2D+vIa+TA0aaquo+b5RqwCZaEQpGmpUchbP13KSS/ptARLOgsNibV+gaFluOLAbsssgejTWBs
nxBYzhx8fOv4XD5IvHjW//5HAzIMDNmBvUJSEqKWiRl9Rixpu9G2m8yaEsHolq82f7V8EfGSDHNE
1xBKN17ZO6jpGXgq2P2SIuIXWMWImSBu/ErYpA6X9dWm9UZH/MSWE8Dtc+uNn/DnCBefZAlef7gC
iNiP2uBO048NxMAX5V+1/B8L6ikbcNvjZ4uvHtecIyGcYuPdEkksOhu+IoByQoJmukqm2qW06uyb
By7QKoLDzn6NzRTDBg0IyY9jaVC/MZpCaJEQ2OKeO3ZGFSBvf2OqJtbZdzekBUn9zUi9YY3BqQCe
TpdV0wLe9J+3fX7jHf4HdnZoO4coLinBx99Iffyt0gSOii7OGvtqLGx1cPHifcZPggLg8X6Pko22
rMtcoyqwEU/81GY6pHu/pluDD4AfphQgSl3sFKY7Hird2p5ePN7HuTrb7ZNQxMEgBSIXNVCdzvpf
ONbARmrdgDJwH9k61fw7zMIcFlUJWxvVE+yPVEhK/q7ASGxr5fgV504DdgozwVX/MxY6zMPptH6D
grYdMVD5kzsIUdyrj7rjcc0q4VPu+mD6zLBLjVznmpJlxj8WiSfcCIjsH8GkzrU6yqUFGkpLmGMP
A8v5Y0eot9D9Wu0r7yW8PvCaEK2clv+iEmDmewgotqjY+I6/l0k8Gb84UdENzF0sdBfVDXQGVyMM
Zl/SirUFc9+qjljhVrd/BrxJUp5fyiz+gLx/MiSWAVHoAnIRq+05B2Vdu2FNY1x7t6sujEE3f3bb
ntz7VV/wDwzRwgCI199AB/3VnPVxdGH/1jw1Ge8m3Pz8Df4VyChuOyJSkiVd7KCNZOta5zQGOPPb
H7CTXhFKUIa4R/fUihj5tUAiD9S/0rofUgYN5TDBQzb/EubM5t0HEOAo0UiRohNehsmBJExDatlP
Z32n1FTqKSIbsiOmmYmU+CCCM3iIVjGj5nOllII5iRlxe0gKTO3pMLWOx1JBJuQVq/O6LVMWC8Oj
iLlNw1V/UD8A0vECdXfE+JgQLnlB2xAsNfsGZAOHrEuLtDqhrWNslg5lNBDPw5JesD3fph7Juj0o
t3+ouelbXrkwQEXBu2Vx4g0EQwgBQzwzQWGor7zq18YXYwLrB9k0MEpk7R03Q2hp8ppKsdVCZCAA
At2SWNKzANZfbmAqcqeFOqCwFPeyt7XxGggEG0LvyghEwgwjC4XRIgcRcpv+qABhQVwYY1mhZ+Za
VzIDEs2R5LGnZT5zLxZ6mq4j7Ti5vRB/fC6c4uKwtCu8FbqgybFNe2r7+JBNai7atMOHN8GYSz4p
DLCkfMi3+X9RQMhHsxOOoJKzc9l8PAi7x+zo7N6nvAsAQ73cuS0Rd9HfDq6oRyP8ZsmgLsW2Spb6
uxK2v/3yjrhdSsmDfQPCUhzFYy5Zv1netvwEwLV4+Wn9XwyVX8XXq3Nhvjk5k0wKbZL1D7h/9UaE
yd88H5rj2oB+9CfyvBJ0kZ6bQsexCNihxvBhz0gWlZGHD1ueXEtWcjoZESL2lU6VS0mp45oePURQ
2pUp8JWxmcspWzRmYEEMj7RMB3Be0TZQZ1IsTRFVjCfAYqMDf+t/SmhTBpKstPpvDAOK7Ptar0JE
Byvvc/H6ZNCPXr4CJAQjCh05WIylihm6ZrSHAGIs35Z2nKyfO6HGrT1KFI2ufaJkSD0qYJIn9B2d
6KFIXmAhsQF0KsWGybRNEbPTLbgIAeWgD3W2ujtA4knrQzYLZFn0EqhvmvndqUdpMkfqpAg6k+8V
mKL+KKWWQ8eMS8BKGIJ6mQ6vylRwOaCSnt6DZLa4OAjS/D+UFSGjSkeZq6PjnJGTExKweyeu70W0
5G6eJ4Ab4XV6krdL24ynd0CgeuSqu2uYzGAT8nxkBcUxcJWpU4L2cdnSYWBUZkaixe6au/R3VLCv
azqXVCcbPfxOnuTrwuVF5Db4APyATZalwfW4uuzE645vRYu3kWEb8PIsTsPAGIUyQA1DDZnfc0dA
zRmPFA4ObC/nxwrgrak5DNFW8LRe0OYEJnQjxSvsDQL1Hr6yhPI0c58JzQNrq4/ttHl9u9cRXa9K
UFHuLXdyZIzuVJ0x6zowDgXTexpJ/gx2g+nAjgPf1xhiT2Nz9FJQIM3i3vfkY/Zomw7Rp/XJ7ixp
ky+f2197Tu5hSdTRfgea1xv/tlTnp9R6xKdnnR2dzfZmtUdEngd3jmcbc7vv4TAYzxmo6NLZK0oU
aL5Nb7ebR/DS1RsfQLAyYIcVQ4n+Td8y1P6b9u8KhlHiyy5mUCAG6SFQvQPZf35FhMI1mj/DzUjT
h83riEf6SIXtMG9e+g35R3qpsauZOlEVwOkXQS5rdbLwXAA4R7sA7Hre6I6YQz5/7cNCGLfSroqQ
vgs2qhh3jheMgg1oQG9zg3EWRpNFyaMTHPp1cmemghHGNSMQKGKXLgz8indogB5DM/+HIBCXVu4q
BKZAWo4ghoekgNhyUHFdkUi0vV7vGmxafncehN1jJLTri0a03LAjx045ImUJE8KKjJUw0t9BWCXA
bzujp0AxMMg31DP8b0CBBRpQ90MoYySpvtCGQGiiozvWnIMTW5hF2AnOv1BKrZ39kLCCGPdTEehh
OjsySe5jnIuZ7GPU0QRU3Dv7amZi3v2nXMgGloEg8rjCJiYG0bFcIfbjr6KrkT9oZ/WfoG4jkqQO
Q97Rn9vZiKNvDyxFYPtkMgU47eG08c947CiiQWLJJLULt7DCcRGfU+UWLc32AP3XeesmOTnRVdtf
NDhZMV4l6ewGZT8Z3ZqsaWFvqx+WTOXUYFRnSdUC3JcLOweJHac3NTsomGIV+WLJH01sViG/yBGJ
1Rim0YvWLFrOKdfTeGq4o0ImyYUXeu422WXSN/sM8ush+Z51QD+lSXUz18SZP29BJXxxWmXlR7uH
KQyviCwr8IYmwzveUBFlUobXYpcbg7nDhNQLc45YuD5syTeBRc8jB6fdgzDOGpwbdyNZPNvbMvm/
Fr9Gw4fKKi2prA7tSgtbeZfTdQSW+aQeGIIVB44g7J3mvsyoG6FHepTXdiijE1UcR30cX9RAmu8W
KN+Kz+XH5D+cUHflBfAHxNKQPUMCP4JFzRTJ1MPrXj9AUqoSj0Ew3q0nSmuNsuOQ+DLH0VrtCqjb
QvefrsQUQTPM9Zvz2Ux7LxN9W7t8m3pwrdtL8mC+ju7k6QDazLtYo8qaa00wh4VZPlrtOPVjZc3I
igVaFON56K0DCxcSeBL038mKsSIpS9jCSVmYKc8ic7P8oIvcoB+07Z39nq9mGBETLe5PwTS2PXFd
Td1t5RkQPNuToIqgdBrspjocQYS+hBhtibnMuMi2yYNCxwPwdfm2nzQ1PjN7oAYHzo3L/xIVgvHi
gdTcugNv8+SwKxiEM2HiaUSt8uNrrVfeV38POKifhVxskTvmpYSdRK08/JoaTLlIngw76/6yUq2G
sI89InhKKpVF+LBiZd6muuO3J5rpUCNBgVmNQbeMPg9J5JqdN8kYKc8NPveYWNB4zFUAPbS6vAW/
LRi/uC7IgPSlIA5XqTz0AKyoq54lT+hP31TXAFitk9Osa8+RDx1vZ7dI/OcHC1cT6a5h+NjtBRmY
fvwDSbEteUyk1g0m/IbF0AXGxPAouCeeb/+dK1chYXAZFmuQHOInY2UusYUyFOwim8fNXJSwwgI6
33F8R41A07tou4sdnkuHWqEVw6vObUEEqJBuPN3AikjEX8Q4uZhyN2m/szFwLLxRrIKB1Od9RgFI
iee80kWsLk2cocbgxT/xOHMN2a7Cu4Ig5VFGSQ5gXbmAwMLXq0/7MlAO9Xv2pre6hqs92Nd1/QI3
7ksjDDb7U+zH/O0G17WVvC/61LpDWYtDAapXs+BCvn3t+/8KyHwcsCPbzqdKLub+hqETh28gGPaI
QeC8gkeZWClF1SicEn5p/vI2p+PC+Gne7TArCmR6zCeBpeq0E8D+yBTVX3Fg6aITYiNR848bcJ7y
6VRr5ZHx/6H8iOVz35MoOfhkxEqic+/JwHRx29cTZpzlug0EN4zi097OuR4A1PoH+2V5EScNX1rs
slXyZ379tehpL5ED647dLIizSTm6Mz9oYLuD95Z58zNf/nlg2l1bI6Q48W4Z4RP9Hl474/zK8nhP
fX4RtmtksrRixCRSyaXM23RxZ4oAqFxNS7kLeboRT6vh0ODxqay3OGEbZxrIYJofyuJPLF8bkrdU
QibSfMBzpY4NCdEmanxEq3N/Wv3lFXD5/VEdpCHdojWhheZXtDd4pa7PYmWQ41dK4raQAkHtqF2x
JuWGmnzwMnJoKOP1FzZzKd4bxfpUc28tbMRb+TIQostdTLEqXINMlIpECoOqW1ECVmixwcy6xH3I
aBzaC0/AzuFBB7qeSOeyrPVxdJ96bF+u6mk+fCKjo+A4zxHwDJv8cHKfWbBWzhJQPcX4lnmWTgOi
d0EeJt0mNvWw7DRYQ9UqBHjqMZ+Rtvhxt1hWKyYDX6bWi3IwkQ+W3BxJhRnYZ80yq1vU0Z8emGpS
NzEbBjYFi3v08kTuksFcXil2uUd29DTq8SUFzo5f9P9omPCYXObJyAwUsd9wx1BGJxq7vc6HkxgP
1JiMxt2pkR84JrH3JrJBFqtMK8k3N7pvg6taFdqBIYLu5dHhtcrzGESSaMgOcc1crR1/cWQdoG0Y
CJgULctVJGViajdPPZwS32vQhx7NKkisFZR2iSp5mqFJqQatsfUilWueoum2b5knqBFcXjlolxIy
l2yj/hUQXhueIA0EK4KpRbSni5XrS2EiW168X04/AZ6arhRgP2dHGTEom79r7txxS2+9XHOhe4vw
oBwyZ5E+7N/grYH9smkDwrqfduWRr3vtPabmkEqiP674gZt5na7Bghzi7pLt7oiIrq1sLl3B8FB6
BsLe7KSpZRWeWVrP5fxCCV1dGdMZ1On/USh5Dv4Jd/o0nrbiwMCBvLNekVoIS9WPlT9ARXcyFFBw
uBTngmgijKICCkg57zdqrpAh0yel/jiIfStZbqbjC4Ceu+miydu5DhP6zcKxtaKzy7mYi/yxgack
Drb0tsFX5gUZ/graGU+tWZIVEs15weRyAe8rLunIppfO6WS3W24AFvx+b1Q49pvKhqarS60XNAIF
MAP9JrkPFnVvHX4decLpxrsP+sHVbrV3/H6sfrxUQLmtbuoejzuDU6krxuTKh7imPeoymPPTVsKV
S4vZE2HHXXAEd8FOuVTAJbxwTV+eMzAsexu2Rjn94SdtN+sF31fawnd+A33NphJQHz/fQ7g4/MnD
2dPEGiJpad+EwgrnJtKOegKJSkJwuJ3u/pSnzTK6DdFjrd6mqZth+fXYEQlzkSZ5BlpMkgvfZjqF
NAcR57tz+gSfokDF/rQa1lHZ4mWf0x0vFiu0IgoxfWvMHVZPSMXaBKMg1k7cf2jeFM5lWlBlKtDv
v50O/I2apz7xQKBEV4iP0tR4vi+P/JSiTvIcKAU9CRII8nTveLi6ACmrR4YDwrhZuWtyuTAXB+Uf
6bZXQ8dpN15Wf0n1pxS148TRu5BLJbtx19bGqw3vAoX3cisAqW/tlvdrISEOPBNwC+6BANJlLD8T
5qNV3Ft2wfzJqALbR3kMsLfco5s100t5SoUbWGM2euzDf5CCq7cKSmwRKjyyqmEYYhs3KYVIdSLu
4d77F4huda+8cP/Z4ZkRLBStl+zV+Qjsuk5Kl3BuJ0kRO/AYMg9AVr0+GizvFIQsRi7tqp942Db5
M1doloIr9PJapwYahyz44QpjWQf35Ct6bnGvr0Npn5aDJJ83PaKF9hsHORPkUbyzKMUrZZz2m2qm
c0ltEAJK4mXKWTHH/0db3mVKcrpsn7NQ2dWIrJe6aVZYI0xOdo9z5cvxP5FMfh9m5UyHiT5G+ohg
9A/1hHXdZ+G9e28Y0zrVnl6GHywtd4NKqzI2QSeMqkrqggrVlinGw0dIBbAhYvVqHdu9lgs7xmY/
xuCYunib6YtQ4tWv4hAuDj2ZJ8UN2O3qOBlNX8kwomiPIRgLo4DW172HCiW34Yeio9OvERam1san
2/7zuV+z1zzOgzXVPtWQydsKdUEvT4I+M4pKkp6YiAfZzdsU0FRXd6BK0+rbNsEjT5ORIcv8Cs4y
HN+4NUt1nmevCvXSwk3GxqlUU36b5IFPwum/6uggZraZ+JFPAg6XhYNDlJd3RL4wpV9UCGcZYt+8
4b6N01d8yOqOaBp8ye6DsN0L8+CtuEojPz1Ww3u3RlIVqGfc82TDf+kd4TaGT5mO7Y4+ETha3ala
ckLN2tUFmm2Dvb5yXYWT+Pf9KAzetLws6gcJy2oNpfOyBwl30iCNgi17dMJywTKQGSxWgg9Dz0w6
nEQeREwVaZUIophtK42r2DdRszIGqZmnAM73/1WXl7+eyOv6kgX9WguBfTAdqLByPIPvPbhSrB5h
rGqKVtYjmRGNC96XLi6bSbT99Bg0P92SZ2vwMKhxvl3fhiSNU6vr8oZ4++D2rFY2520bGVtSInoW
FRwTe/ORmUcsn8sMSWBnUIyeFXsECzmO38yt380X2dKt7u9Z2buNdZFJHwH5dTWP0WgZ2FLP9M73
A4Ob6ATcgD+CoLJbMLRB2a4vIw4elZCPiEC2ORx/Sv/zCJXCG6zNage3SuUM3oXCsrRRhUPiGPiv
V67mE+05asd/8SkQOXO31pq8kW5Torpf8KCx/xmi7JSotj1NS92Jve8VuNVkVsY2pN+7WH50shDW
hSmwdzoJK7BxdiMSgW58JNWMW5hsdrdIuUEV3dth2qHrJd/mdnRI5iBOQF9JEEr+aX89YpUvf+qe
P2U5ZaY0gtVUswsHLj8+B6u0ygu/px6tIfYftsNStsU+jfXHnHludfRtL5lVdiKVoV4RtJdq3Xc3
VSOaASoSkc6mh2pfQcvbxhLSZlyoNhtlgBpQ8gBgD2c7qoAgpCtPGIrxttu9EL3kxre4zUO9EbZJ
8OHOWCMbzeDgoVfcKqIEmyplGnxpYqI7yDXDxAmr+HUjog23EmcGqqXnoohZ551mPKoOQdXtTp2H
r+ct8dD4Pnf7IweJM1R1UFcp2PJYyhVL7fAm0U9DCbIKpa83NcT4XOZlDvIXRvwJ6/sVqjcOKiQ5
Fl7zpUqIjN1AWYiIs8HwO/UGILW+wGqHwIM7wfLCcEtkLHLkOej4CTO27seB9j4+xiPLzf+3tDN1
ZfY7bgRtT/W47YmmW0qDJ5HDsGeLUd7rFvUtoH9YPKxAtIa83w24NqIdpci0K6PJTvt16ln9YMVh
MmdbMKJQ5k4gQI5HmGeCgs78ogoX/QqYPKW2g2So1xdSxmo21r11EdyetGK/C6RGVMMeDL6MLJkd
mMrR+1zMnGQU9cvzgE73U5SvW/xYjnf0MMuLb17SHcgmLPpo0OZCEO1xTOc1KdQNm3hiRNLFSAhQ
vj/STB9IuuGlsF4AmWhVdmiES6egHZZmPaNePqKp/iF5mDoJH9QSyGkwXAJDAkC0L6Oh5Fm0pIaU
YmsTkU827fYG5mEsa1BjjWsSgMJBCJYGU2LcjAqc64evtt9V4Ys2e5ooXudJIqSVL521rZ5XbNXW
5ZTRiijYbJD6ouIQVivqFRGTKJZK/q7fMaVGI8S0xZE85VvuFO8PsC6AQaQyXrGVEzhw3O2fSXeY
FmsmBWJMKOgWZqWwT8Ypg0r8AN1tek8vC9dtDJv/1omlkcv0pazy5dzbSdCOrz0klZQx5NBgZR3Y
Q+FqmN2cHJdQusXZ7qfe/k7BroztyaqvEqmFIAjQldQsgz2yndzWd6N6C+c0K3qp5BosQYMAyxAM
FZLHZqrcdVTOaz98/4a4AO+pRIOfbnqhuKnOQ7oTZVGlYDVT1AzIu+gyeujkjSOgSCL3KsAmbe5t
jHVoZNlnP/xmJVGkSXkZGQLaGyPC/RfVhSvX3irkTHrxqzE07tmYC26QhRcZGq1JqiQvhTBq1yjo
tM5qbJKHU15uonsiI/RzpW4/LEHtO97qp35mHu80EMpfP9hFj+8WyrejG8giFe65fyLxoQPtuyLc
PmFtQ0drh5Lnzc7q29bcAJBkf7Hj9qqkDXNMR9yr1Ece5gccSkd7UyMxzag90gd8zSsxPSE9vo5N
COwnjxd9K6f1jjEz8l+Tj1g79Ft2tbT+DmPxM2XdhViI/8yhV+WKArZ4AzsUL4W2XapmmfWkNV5w
v656WcOh9sjpddn/etJcWTzcRKzBHt2IccgMX6ClyLrWeYbP+r3Fw0KFUDtfq/7P2xQd6Z4E+Nzc
g5JH781gbDp6VoyrIWWQ5VnAj2lnbaZqskBUVYRpgt/edBCJhV+MvRgTeIbhOOr4DSexrhXdUpkg
ku4UBECYG9u3/oeBSd76f6RCMiFBOCbhycQYHKQHApyR34ZUSvapan91WNgR8wInMNGBYRLmX3Ye
Vj/ElnJMAYae0vqIYQGdZwKBk/xX3WslVFnUQmEARX2lF5vlCxQ269Mm9mBnGGu6VgwjcyZ5m3N8
eGj+860wDl1uojJAI2efV60NF+MlszEfLHeKTEEq956kWfII8ekszEZ0pg30Bc+woZotRmcyZ6mz
6Hvv4oaEUAMa71cd7fOA73c0JTVQa9zbFQCrA6XBoMZ8545AasWnTTAldlBcHfV8VTOG5Ai6Sxu3
/FqAPzZItvQLj4QdRX9JEOaBWkReR0vP1rq3mbWdR5WS4SPa+esbAiZG1PLg2LEMvuXPCijBCOki
0npwqi+NhMb3Kt4SlowvRslP6Ht1R/0PUsqAKph8Ce5NNlOauxYyQXPxWAlz2i5qNVsHEIE5fvfQ
ispK73fd2XnIX8LBp5xMmm7qAdY2caxkQAty0ECSKfaWdxzPu194yvg40gpNGfUZmCh/iIk+9bU2
dlvUkk+jWd9AlLXCR5NmiNn4hRw0XFKuVjWLIgqLWSFwfCJ+4FZSp1o5gbFXTW+leShgAAXkafn7
G5XxgPnX7+nioVPQ1hfWT3TZqvNhYTx5L/Hus+rBlsBCiEJObM0pH5sBxFUwSectj/Lm8qqPA0uO
9ZLbZOVRHr0VukC6I4k8jIUCLW0xh6RaW1SwmLmZ27Tnd1zHKEzrlX3KfsJ9d7zBR4qg6slLVc5U
6GQF13oxFZwMaOF+GJaHCFe7gdcL8Fy7wKmkgjOQ6C8zG0+WfOR4IOZk6lbGPOVvZpVCPQsEqNqV
hMSnUpSCRCYPhPyLhsTNNGlAwy5jfYEmtRlcrpuQmpV9mxbXHMAMN4v/g2ZBIRa6tQWkQaJgQRfU
qYtzBz7Yt7i8NEY5oWOrCODYKuPOaQqFxPxjMVE6CyZR6LpDxW1VC0ED0N7Gjuu9hxMPDNmBAA5L
56PZNlPqwrgQai85Xht68WfuLhBC1pFMjdSNrKIna/QHqWzdZB35i7D0ZMbUNXIRybkYxrFgTpwc
ccPKrVWVftbHTSbFPknp+6coivGy0NksnIVbFGlhdm3WlqY6hMSlvuJ76oI5u1PpGPcONWOQtIaj
xuI7dU/Kz8SrV7zrneM283isER+dQLTe3dhFNlJJFd/LjBk8K6gq4VBz2pcTjrpEj2TfyKMl/cax
SMTRjnaIWIm9q7IFzMHhKj9FVUfpEWF1rVQWzPkpsSKKnZTOzc8IneSMPbfoVikqHMfKFVwgCw7i
N/LWMj0F44dHzoM3A0yduh6XenQ1JKJCiPNa+qUtMowvEVpp3dz/gsY00pVOhu6yle/zr8NDObpu
FqgYFTB12ykLcjmpzOvLoP4Yek4miu/17N+17GomBLTxQQFjMe6N7wNE69eqF+H0iOeCfr7qNNTv
fSKORg6gc6bz1N6BMQKrYWVvmbsJQYnOP+ZLLp5jYEWunG3UuPchFEfhnoZV6MS5MZbHfVuFrV3W
MstY0jIEYZXw+P2phckxX1bOyuiTGONXcEgjQ/64Lp9k//1/PSSkWwwgWEitWuuRt+8qTooPIDF1
t71F0OacWCpLswDNd9dgMYRGMHYsBVDNrH+PEhpbHxwNkpFmkEk3CmH89T3El//f3IoaMzr4CrnS
WD/t9qNoNMlOh3+DPk0JkgmtQqSOunz3lyXxy9LJ4pcZvWxhyOwin61tluDACxNfXefJv53+S3RK
Wh0CakUVUO6X7CTX/OKzAKkbQB3ugzhLIBkvuXWSJWBRem8qLDzKlQ12r5iSJkrRrP6frLHf4wLm
bLWJQAkpPoRGeJlL0DiiVyj7DngBJxlTC8Dp4FbVlET6y+FMTSx/FxIwuVXUzUh9IEEyWkpESiG2
xzT8zTDdBRh8eu8a4Q6cKtD+mlA1GV1qmFwzFYHSU40XuZNyJeEKdujkI+lKZwO//ZX1Omy4pU9H
8CmxwlQ6/WIFneM7usFlM7ChpBqbiSryUtg1yEz3iTTK68pBKg6QtHJwbsPJcsT4ZUzYFWztwAim
b28js8Fmly1AXND1rtR0bpZvLC7sh7wJpYZcZG7LNeMI97DW6g56RUehauQKCwsyCvJxExEOW3lF
GS0Ac98RLxjAafeDJ/vBl7TudbnnQQOO67EVJ0n9gY+FmJidQ1/N0rY/ebJBDeT+GWrXZDRcmk/T
xnlfpaPAVdlSOTqmGRsH4OJhBOUXkrVF5TtpQKcSZVCh8OIAPh1y8/ENyju/14NGaMrhUoipLair
Z7JoiBd0WMkVvW7wzny+AzF8RkaLg+meDdy8zTcAHFMW73LVCKRTaSOAGUe5/DYIiaWWh7q18bWF
+JdnMtVnbIVGFKI2P+/LVOKkPGQKY6ykqDtFN2t2CBYEEZDx+tiQyw2/GnlEqMPERF12iYjq9PPl
o+bKxAw4VTpAgJeB9L081+G2fyzL2zPnX4e4B2oFiFQIea52SUbCOPrO4EP7d6qqkdRN9laKQAVZ
FpDBakjBkifj2YKiC0O3gk5U7OAZYhDm1Bq5PA9JhLtpznGaERwIhWeGO+TIEWv1CcFowvbuUzlr
cyUjYwFP+MJtPQf75IUC2QFLt6doZSNFDEdMbmt/MieauBe4WscqfGoZUeCe6ssqi8FMcE8061/r
HxuXRAsFoAr1Ma/s27AS9qvEigXNcsxSF2PCWPbtDR+yvJgseMv9maPM5N75vFacJxYPSCPmm9CI
6MQJSe6/TnpqlaRFn1VwjFRY+34XQz2OS8kvMMtYZRz/b2ent5+KxL8RZ1usayyNoKq5X5Vo4LmP
2g0qRR1tX2mRvg2Mun8GUBQzLUQI6RgPIgZRNtdOLQ3+d3W2Oyoeu1lEDjiRqvnS9Op14zNxOL4Q
1sWwn1OqKwLBytcobq3h9h6iy505QeGPdjFi5WjwrD1Wf8uVrpuSQrUcqknbxgaZonLnxUFvMvZT
zPjmbhczcecRebnd2wMJXuuKE54zP3Ezzg7tf0mNFAdb2cHCRMiMYCS8/imaONz3QLr3l0ybRa71
eZg3z2GciNaYpLuZuEgW4ZpDeSlVQ7wbdlfPNDO9lfxXI/zs18KUjPRBWiOwBE6B7i5yNY3iHU1m
ZgYPu86G3Oxd/cAf+846tYO6jJXAJPB0tQ1jzUpGezsQuwI8CssF50XoD9j//y3XS2kRpED5lR+o
Hp07sSb/jCDZHKnaTlLOzUwWecYCASsUnROQM+NDSzWLkf7cgqkVwT6PQa3JjO38zjjff6uLvPRs
IJQdKoxYRWXJw7Bw9DOOX9QDrmQBT1yctm12RY5uQty6/285eBizSa7UyaMfLVm1I1XY6WcEOMMR
lQ8SARI8RMnFB8HiSGi30IXLDo/o9VpKYNZly/5fjy5JPc12gnqm+0TabAJwuwlcaEXSE/4/2NYN
g3xqqOwgt6sRizpwQQcdG/r6v7L7XQYOwRVFrw9gpTnvVNI0+JxiXStB2BMY6cSFtfnbjMYpmuYB
d5B1mct400agbjofVbZOlJgPcMOfH9D+HaVPejQCKGtZ13vplhnyjIEjuWVeS71e5BMJwZ1Yxd27
Wl9Yyl+KIl8AXJMyYt/oe68+v6jvlCUZyc2zRCqhf8WjkabLhP0DPkVx7iJJ/WH2TnKgNkwR6Bmt
U9jn2YXOgLjinurhCaEPIoL0yfgrQ5WLNVUrrS7jQGTP+8qbUho7+oTs8XAZTevIsjJfaDEoCVKz
dMUSbekSs9jOB4Im5mvmQMSDwnwqah+BSb7RgU/dm28CdjxRy0Wi31g1aIwUbfupPhfBrcIYIMGc
wwWRiP0xvvFuGuoJQuYa65V8u7G6ZeDpHJ9p+SWH60P6vtlh+swghet3vArdc7TZOmk4zl5vNmlT
daaxXD9ue5HI4V+42sB6G8KDFFHy+s/ATMoTg0dFTNV+DuvHkByKGdlmi8mMCAm1v+q0tAK4cmEV
ek2Oz7/n6+9k4SIoxC1EftWQkeL6rYJtgfBWcwnsTNoEe9Yc1G7zlGTbkMvrP1+zl+2BvMTc2UvE
goBnamaBiUdyx+ruqcMFXuFBMFwR/Y/h5wSUurRQ+/2dtC2g9+FwTmupaXdhIUFTiptaJSjmFw7h
RFZYmGZhxXrLqpgxcfgaCsA3O0EczDVVW6PikQ6Yv5Fi4y1ZpcI/waa/RTHHNzKMN7Nh65HRWOhG
t8judoxqkkNjsnScQ0cH4PdODA68mHAAUrgd69xUS6bnQD7HZ7CVKpWKyJ65e4vOS/O8w75jhjjD
XK00tnHY7QkGQcAWOwn6se29VFRZB8UvQPdtGB0+TqghF/c3nmFmVLZzTW3otJeJxsIRXPkJW6jF
AVsTBCV+UV3kmU6HKFh7bOGg+qDeyBqGGuHsNAuQaoTq5U5vMfGMQCzVosWHLlkLwUvlZ6esf6oe
QPdaEYbjFdbwgsbZL1fLt9GzDVP1oBfExt3dV9uMARFbyks2EQqCor1C/5uoBJiT5C5KoclTXoXt
iYlepms7Vh1K4SimIKcYADjyNgHXqo3Igcgs+Wvwg6ei4IzpamoNExNiQufoUDgwGsOq9LAOXm1b
HpInbwabwXE2UIKgEif7d4ROmw9DBfrCGRzL1rCj4BxcBp3OvfGg49tAuulgwyDw760x1LEya7Gn
oCwXThq6dqQYx9P58hJIvNWOMApubXk5JZ9N1wsMLQC3zz35a9JosMtQculEmPa8AfinBQ3nRsNC
z+t8WdcWAKXKjW1QaJf3YDykt7Wv/KUhK+7f4iQqH+9QGz9mt2m8QQvLIZ074o3n32TKqEPauAc0
x8PcJapK8w5y4kO1LfWdWlRGIxfk9+NY3sknGICT78GFuzuFGwJt+C49eKx+8g/Xw3l2EmhCWld2
5cGR9EgSiJ36ydD+2rvX0CAyvDcN7mxTSQdj6GPKJfrz4+T4VAbZ7Vmo1s5scgdlAxmYZejfHyLE
3HZXaQsWX1wxcyHx6l4n+C40aH80b/DfEWvymt9a9q6hPK6iqDhZ6hNAd4LsXyDj2QtZ2XtgUkde
rjMFyt2Bw/IT/t+z6jC8VO7xNhtj1HBuw/QTY5yn6OnqqhFiktDs5aiff8qjbzSyLGBk3fKjuyha
f/h9k0BSFwNfAWnD6iX6t+6p/7UCaukE++La0FPTsSNR61Aq+HcN2VgQ9L87kiTx8wz4nrgPwqDB
RHM2EYB+/MrkBlfuxb+AQRqDxWTkcBfooLol0EywNwbTQwEXMI/Cpm7ubBnrOuF5qI+LRxt6RWWe
r//hRVLUhM7MdcfifBXZurFCNhDrK0fti3E4fyA9zkNmkON05wMV7kykx47zufgo9Yuc/+otP3J1
kmNwmdK+u6FpKb+8njcgYV6zyUFqPTXF1Urpft7QKjDxsnsdPGTUWqcx+asZZpaYVOZGm1rPtmeP
4DNL8m+TtZ4X7b3IOzIhEw9EZc9vF9O+WiJP/4qyb0FIjQkepaRmfSkI/+x++t7hfj5cho4fgW1L
UkNI07KG9R7WACFK+1vESa0bEBNilu86QLtK9u109egmQq1Vmz6UbiyrwcJq7wLTDpo8Twp+cA2Y
sWzSbyoYWUeUIUnGQ0B+SMVLaPfT9LoKUcq8l8IxT/LUZUKJXPLHpZNVhbLxlUxc5E9D711l7UyL
WBgulzVEN4zfMgHHgjOibLs4R2P9FQgK+pcyUIvBHshUeOTdpQiRZAGc1r0rN/RTC5Z7V2zphui0
EImYGXpLLkBrfwvuaK2+/NTOLw0UiHA9ufOR1SrnqXhoXp2R4zm/+tIuBSwZwOeXi1MEuKoG+pRI
fEVCnUiv7xXvkc8ll9MdFsX6PrPfX+kUjdCS9Dt+Ui/cp7FSiwVnmWcs1s/SpODUCY/4HDfqxLJQ
4nWSsQzTlHFGJyphkJpjtTohWrDjRX9yUjdp34+kiYsvxkLSrCwtKFnrQFyVewuujC8UYDDmLun4
ZLoQisHTzUjfgp7Ls+hyGnjFG33mBBvbZCWfR0kCiuZaxwMp98++oTpMvA5TpAIHsmZol3UiUCFB
QYt1WtSKPhUqfCuC6Iljt3tfrdznhxresLVljfnpiG6KJxmApPPqysr86JYf6k/Znooz+r4w+zX1
B51P0UCajy21/8VA6tvNltR4jxR/JN12pTB+EAsG8SU+XlAFHlcfOqrnHgYiZ7QodGC0JzsU57o9
rH+1/L7nNeF6yDHBI6db95/YgZso8/DPYHeL0vaMX015wvm1yji4uY39I8SX8t/QSuIvVrYqmjJ/
Fw2CMR7um8sCuxvclAkSjh61jb0X+cC/7fYYbdLwJEEWYji74dO51I5dmGogGe1pSkgKJcHT8nsD
3Ie0wA4uEphQ1mW9SOGNwTtJjwGklWvj7iDmkcsFdHjYyy+Jo9CyzOvXDZUARsaQHeR81L+5qFOQ
MfXNqi837SY2Ud0RJL5hye3nFZ0A0MC/eghk6m3+cLYk9044MFurMaEeeNaRXuoj5+dEqITDM7xD
C91SzBQSPkbqPhd+xXqlz/6+bMncaB8zUeGhLDnc3uzFz+uqxWVKHlGHRLPO955fh6adQnJNq+4i
79uPSgv4oykKcfU044XsxIzCWltHYQptCpW552r2up7L19HmGS9jFnzK8dGGjlSJie/p84qqReSS
VIjD/Q1vEoCBPPL2/xsnxNL3c1WxGnVCAZz7nhbkfVMKyIscpiw9YTIEPyuL4MCqHDP+hcVsLG+1
q5QEBvwwocRnTlsCNMemF3uNdEWinNZcvHu9b/tGB47+8H1GNWECmFR+r9nqDzfCMgtnl9CEJF0b
6RUVUAy+AkoPFbiA3z8bA5gfbyYzX+sIhbIMOmXsP4xKOko2StxEhm0IDDnznjXfDndK6Ha0v4e3
Eb8JWXNeupYwoYQ/9pY0w07DA5DV/qNJI7FbsvTx+q5r/82KAThh3ZDZjjKeuBhtzcCkd4Edm9hH
sg1nDgxk+w5bqnxzpym/5ww2YTT3tYrBVzb7lqvnB8a+9fACTl2Sj3DCoWtwVxEBlbcnRCNpghlJ
ZEZupOeAqL34KrIzFuFLPV3xG3oY+QAUPRjEP3ggTAJKlXCuViYLaNRpGeduiOjNIdjsvdWYSpqZ
QeStmEEgiUtOt3siltn/VpquqfVZdayb9kA3P7izOtuMr4vfLqqzIfSK15Lk5m7A6jlDKJv8q50i
evMGZd3KUc+sJaf40OeDRJ5wa7DqEz2sXdFz04cfOc8wUj1ssTX85sxRvVDlxr4uC2X2ui1kLOzy
P8el7QR5aRkvQ463chA32FY9CN+oyfCBU7ZvSf1GdFyADb8ipI78B4eKZ2XOsIYiBygV4eCJzsle
KoGzVLQjOgISA8gJ/Shg1WPcAePwSGFFR/B4PQhgft30+AT3T8oC91iM/kfciMPU7Z7Gachwo7hN
xk9LgCcu21drixI5qFc13090ig2ssb9W/274dJAPY97bUlcxEHFBnEMSoIOrs6syzaZxBO4VmBH5
3iljZAB3OdFv3H8NqoGPBKP65/algabkuiXX0P+66+BEDEuY8MpWP81VCYkxYLLKxRED8+83rq6C
PKG6AnlXtZEBubDbNEIUYi9zLFJ5RMYuCgKdpk2nf66658LeulIrHFjUyKAim/1KVtSJxBounDFK
yscUZV9jFIIbJy0erfmRfTUEMMNYFuGfWtwU8H8RhzO2Uu3WCU+8CMP3Eui+Xdkun480eIVWUCec
C9bAmyKuhpofJYJ4zOzsbjJ/+bSOqsEjRY6a9TQlGowo9Mzq8QuuAkkuSvhDP3U04uFOYgtmo4aD
vJecagQOcSAsRKp6M+8KFu7a7ysdql+lvqCqR8Mfedakyjr8I0/4fy2pS9yqCEpHGjZPcz6OPaJx
HGGAy6z2Bso2KL9DXWrEZuPJSfIX1o/H/Zx2CnWXTVyboLXgbMLLmeyfQF2MCIWTIvQnLdPZU5Jd
vuWpAnptrHfrOMewXd4Bzxd55/k+99zSKgb12767XNgRHidFgruwZ16IajJWN9YsK4dJEh9Ry+uQ
6Qz3O60gcf+Xc+EdeVe/erjbQQwUvWt6xHiKbRTTD0j5ZA1+udkmfS+fnww7dPhZIoJXWwAXgmNc
1Xj82fkFc4RBOe80tBgVUbt2L48Qgowm9MCxxW9lXPjDmgISXKG6Yl67rOYbldKjYeQdU3+2Hb4R
6uehwD5r3I0yECVZh765bPrZc/1BsK7Kcq3Qp5b1O0ytEMkETVFXOOA0WSjhOSRLXv6pAW7y7sbZ
ldFxtjCsOMVj1XuU77N80ZPjH9rBYYQwuvjv3+lz2oNC/dJxWwqU60qQ+NHLh/N/LNV3OiUnT+uH
TLVWaS/omTOUQOE+0h9MnhkBhGHdVrNuz1RaGrhMtfFmoeMxWgp5nnfowoqo3ntOV65POjoTcq9f
610yZnoz8pktAMgAeB44Fd3Uaa3P4xJsBHYwfjHGeMsvFEA3q89RjzRR6L7DL1YwqzoJdehgDtDd
nbWm/Cjm+aHdICWMAX2GSP3wg/NCIOZl/twfZE+bnnYbglKWi91zJRNS8feZRA2lDqf6UcfkPvvb
hEaY+2wY+4FPniMre54Gk5e2CEnWkDlregu5REJCb92gKOt0TWieqQ7LjA+FmI/+SQk3WQ5Z2EtP
lND7r6zR35mktwhEpNaVtgwyiQ6rkKx5WeKgZ4vdVoqDOJ1Bka+q58VktxHsbdilvjfNMF0TsyBJ
rj5OKkpJuEqelPyD4mJa5JlAgD7ZCIrnlPO1Y3kPwId8Q5KkEzREWtJOEW5+qLlRvpA/cQZhEId5
XxNvnbEYXR2u0kuxCXIDqW6JFHZ8hiSe14N8uVkdA2oly1koOPmnLeJEtGUPZw0ZIatE0NKoOkVA
lBt8zTK5fBj4uh9HKi37WsDBBjgPLsI/DeUGrhVH74VAZlNu+WAHw1DM7D89XpSzvcC4tYW0BctI
iYCR24NUPis+VPtMP731Q0mNNBVwvab8Z0K8d28Zs9ZBp82n6xvSjxwtIKDzJuXCBiO77pkkjNXG
HLfJj0wuIKtYqiQmO40gZjFUYkQ2rh/yd5n7kHy2xe/yJNLKgwys2t0ml4OC/k05G/QoczoHJmYY
lkhLC+jibWIWfngz9AFsFBK/McO85mTAZ1OBebubBr8sAMCVrx9hgGQZpYG4nEAC+ZBg6zgp7IVF
xmIyn7LpCy+jve1jB8smH7GAFiZfVkmmZOhJx13GrzUjffvIwGoUdNEQP9o0d6I/TyqbNbs1rZ8G
vUiBHlP0P7pw9YYhg/jkWItCXJQn+qvoE5Yi0t+FP773tSc/Difzu+vgc+LZlbPDxKOAYsMluN+A
4NemnpacOo8qdNUK7GwEYLj7VU4JUFrGZ/Ouc+D2FwKo6gCm3F4ROyzFX3CWukLJSQBK2OjYM2la
bNccmXUiVLQHuWRl7019TE9LaXyn0xuAxM0pB5o+DE1Cpxm0HOI2uX2HpMVjGUnBlWQ3KHMcXU0G
RBf68cV9Kj03zX8JHCQrV4MwlZWb6iW1Sfa8k4CcgcuKRj0ZtMAD3tgA9DY/GY8YygWeE4dEgPQE
jCPHenfyqsD98l0c0AoebwrQgXAofjiIMu8rjd0vN5Zwy33UpxsfNBeRWbR1Voq1iT3udTWs6AhO
W5Lhk7AtSi/rLWEw9M+LEM7kjq6UgDlqGdoDtvw8amfE52nz3SQjuCjz24EEjBDrRBdIpyXQXaOu
hNA4qZwGZFYs7TQ//9i67sKfR30u9EbxoS+ow5ZM/q5tFTAyK0orxl9rpBcACXmvNXaVMv7FYxo/
IS02vOUngUHhDb+kDXImG+Mh70cxclQGT3/7o5iZ/fdigYYrdBUaXl/3Xx4FHg+z1cJpGQwFdMCD
1+/xyeY+UYXjpTziYvPRpLLYFiwJSFyOLPUOY+kirDn7DMy7rbKGK4hBxQVDbzrivK65FMwOeo8v
Uu18VM8U/2yeEQwpHdocerm/Z+AfDhgPF9D/iDGjuS681YZOhcZAf+0svCfD2Wv+qVlr+o+sQ0DQ
iVKL2dGSzyeygdbDvyfPcWmgmtFBDj1KkFIKuC4iVNk5iB2qm1EJs/HpjXx5inlMRYsKB3Lj5I2F
5O6Z2X/PFvBUYEeyc70zZGVqWNsJhmO61025dRspA7UheOJ6RVR5cIV7mkaPsJeaTzIVaracJbUB
U4mguAmJVQe990v3+D+NaJGOMLlwCXNXExblbhcLmvMd6GaMm/pEUxTmxxoUy35xcP0UAvLcze/T
5olch5X7hoYEvy6KoZ8gAXA0gORJeQRW0UhAKzGg4BNexVQI0sE/PRVwzoXPE05h3qEOLmRYAPf/
yyOebNzSBsra+rSP1ehOiEujcTJsTVyKxN7crsw6IEWvasD/DqIiwPTNHxy3jtRpSrMzT5+Be9dK
I5yJKy4aoxqs+IFAGjXDokdLyi2bMjBIw4CuPDU+uHpWKkhoxBqDR9skTTxezJ5hZmcBuVAI44BA
Ycmm4YISHwn3Z/idRevQYzyUgMFOxix9NEJb53RTyGDefGJlt0/uQYeEXhDOEoI+XgPqgcKJdNg7
PKrC0DXS2bkynYNWtPAYHcazSFuFhxTwTKsSjkBm63Vp3/uARBsFDliuWVhts0063OlFP6TtMp6j
WGC7y1OBAaeYMjG8B/V3QulknQcnOKaaF/7xQOh3G2/PjmuL9yVyaxgmuqeqimUyOzCwLFzU7KZj
W1CbEqruXI8S5EqwXxrkFSknfUPBtnezrwGN6wwmuZKejgbgm8kEWy6CbL1OpehDLwETKPXLWPZx
ITzXGqdCV510+3gd8z5YVN2QBvtuLkMlnFZXBxEhF9P9fnAy8OgfxE3cTIThvVNk6tJ744rdRVsv
diZi5zViN8WQqXkNnsvf2kSO/8o9X+zo5uW4AtAnhS57q5VD+5egzanc6vtuFlf4V9E7/bWj05We
m1DY3RRsDxr+0QayA2V+w4mc5xWzGLhe4anNr97TXuWTbZgPUJ+KOI7O5mFj1TnlHN9MP/kQP1sF
I5N2xwCQLC930KCnVuVb9DSmiNV0u/WmNc8gmK/Y/s9oXl3QTRktYAbs8YC7DLTnCe+6vlSvdf4k
puO4FY8YNia6udIpgk5sjHa36ZRfrZNmhUMyDycXkAADWHsqKm6Z2Fyq5NMXLIKewzBkv+GMyLXP
w3Nau3N30KsNGfAyqHDbNYHwXRzV49hhXks/W+EzKEVWi5Hwa8pumBnmMwwks7ZYAO1LgWZyuhGK
FunEBcD6DqmEhMlzRLEEqk1cjDuBnT1pG44TuGKBkSnqGcjdRLUSPTssruGIRJHLiypanrr/YO4s
57XgjrY+7g/OvGmcuscX1rPvQQW4Sxp7bs9vcexDxFvZXqA4MFP/4GVR9N/ith2ez20obibpe+2T
LxZ9L1+kkZX7cPmlpmm9/WsuPXJD28G0z2I7Kcvw+PCiAjupdDZQdJIO9p/MHhcwnor7kIxU3piK
1WdGCAwgnS3jgnOUgxVZcwW//xfWtIkg7/EeglCZDr6hAbt1Bj0Gve5sIY65GggdiIo8X34l2cEC
gkiLA+gR8kl45QdwUwAoVsBJ6X5CkKoOzuVBX3wa6Uyn9c7c9/xtEQoxrnzkPsEaRRKqwlgRLRvb
vHm0P0uiEPQTha+UvCJwHJ9CQ560QJTPC30/wOh/lAi47Ua0hn1y4E/K5A0TfHCTRtupoTbPsHZ/
t3hC/ioybRnVLrUt5DECj4EP/pGT9OIKFL0eWjOa7LsGTnDeh+PQj0XYJknFWhqpBmxamKo8DutO
2mW0euEix55uotTW8lfDDD/KjeaocnRWM6SN0tgqY7CKyG0+PHc1niCYjAFxzM7ReH8OTPbSuirl
qys4JcOvSlRM7JncoLabMqPx9X1abOGeroENBHoU4lnRwzAMDOw9b/QCxx7qF7ZFqZ4JE58buV+u
AfCPgxlM8PyaWLzjDbfVmnifo0Thc3hhYDnhPIDwf+6bf+XUEObDFLnIw6hkJ9O569UVwljb+zY7
YEh78mH5Todvb+N5l09vaYnL8zXfpvT/1egu0ThuYBUAoiHzPn8ESnegvHeuNPt4MkzLUFm3sG7S
S9urk/jsuN4sqrTmJ9quWXi7CG7xdEJwxR9+GKlt/Y7xdgH5SGtbxCGGQAKcpvgSoTqZnQXPvr0q
FV35jC0HNSoGV3RtPhgda9O039VaOiXA9FLO2nlF921lssrwxAFxu7TWhRo6rXxJblulrlp6KZ1H
1z8kPmeoHPvxD/I7Ohtl1hM/5C3wxpMr/MJ3QX6byz0/g2t1V6Z+Ype4lsRnva/hMH/LqSZu7mn9
GKEodRAfXQrDBhALm632m66kOD4lsv2PL1OTV6cyBPp2K+bUpvM0YgPumbJ9Bg1CZQUoFevfO8LE
iUeTslD7Zy4ow/++bLpPdLQ0JMMaOqaMS10aMpHBdAc5SR4VKMSO5z5sLiV0IdSY97FyYPbUIHug
sM0aspCb9BdX0isSXeEfMjWPJbCEjmEzJX8WSq06tUrvWGRy+/+cCfc2VSFtvx4njnOSaNs0FWS0
I0OFq/ROblmCCqHfQAE6dIP48/SjZT0HO/tIxLRSp8IV3ZAs47nMN6o/bLKv2/wuvdIbRmVVf+u4
zU5vIcBQzkzgJGjyuAgV4loZazZGLYRkl3fcOof/evB+x5OQJjTlf8ptQiPSrtRb9d/J3DWPMXQg
0roHMljgger7c6dA58IgtzbtNRK0C6WZ4yhV455u+pgy0XkFSlYSX0yMiAi29KkWwiI15joJWh3U
GYSFlBZ8afvcn69U7zclMM9lq2pmRQAm6jIDf0mUkPW/W8qABzm2VBk6ABRdFeBK7XdZn45YhtEt
yREU60OvcWufXUQJSRYrrJNojYIQc8LeYSH3V1HcmAkYFw6JaKfl7pPk0GhAEP2aAzxLzvlKH2Hq
Gza7IEOd1qxEYO8s6zHX6oN6+lBhMcD5RK8/VbZDugP52eSLN7vp5kFUkOQXc31sQP0kIMSeYlZ1
ouay4IFSZeUdLfoDsyBcZd7yTedkQ9jFy5zfRwAtravVHK45i2gaog7Jt9/gXb1Zc8R1Z00CUK5G
W/+KUgeya/2UgRHtCY9Ji7d0x3H/H2IbRMfh1qCysTlOu1z506g8BTI8xWFQqBITO3ZjwscNVJQh
wLwq2rS/8DTMb1MR/4UstyDRRsq2gL5Qlq1idI3ReODWfnX/LlNGlpkKhsNm/OB84hpAt7P4Jl7p
6dHUfhYKxhYiIzVuKEhxR4rwu5faOnPLFq7jI9UCn5oqHSJAYS0PC1LDFNyKGGbDzBa8r58mNXAL
26CWsnv7hzJw4QT+Rfu32nPs61wiFLhaFjQylXNJU5C2GwkN0MKRFwygVR2kYlOxQWCiGhJtIFF9
2xL62PFy5qFp4awArsBE1VUauLSzoAm8FZ7hZ1n8lQ6hJ3ELT6pXg6dzgRVEU46XJLfsk4FP3+ir
N4c7BAo37ZwAIOXCqbDOSVK04RD8m1XsSDU3JyplVQ6S0q7car4YkD0F275f4pGpzOPw6i096zTw
USMa1ThMSFboL0bonorRBcJ1EZ5q8g+TidREbdmSQdmeDHz/9ncxvVeoV4eMNVb5wITTicrUi8uW
ikMCKKXFe+I/SBC58kpRPifLbNB7WPkKppM/H/khbviSeJkZxch7GcqDVs++6incN1/yQCJhp6q1
AQmvHuepJ8orzyKSlpIzclN16fnmgGSnlPHIgELs3GhMeLsoIhG76QNJyJcAp64N/7DGaQvCcjNd
dRdecTKuZLsOJpCrWseJBvqpTx6MPx8w+SjQktI9jzzMOzwZF3v3ieLnEZCa53/i0XQZN4qEQ/XU
ZIR7wWPhGRAUHzyqF18dx5lKak5bC647SuZqRh/068JQA1cNC7nY1lVEtbUeeCG+f5QsK5tCY6Y+
xA2ENHUW0r7Np7NXnpwr1qYd/c+o/XkDbipKBi3r045tSVb5BBWiKjCLJQpTrr8GE+wpxruwYcox
iU46/UoUT4caQzhV5oKvIz8Mj3qeZBxmQ70zfr5KhJH2wEImpQJgo2INN8UMiKJF9yZcOq2NK6Cj
XjAnlTwd0VwiseCObY2T0P0Kq/rfmfUB4YY4H9yzn3FjDMX1NtUtdRw02/YrflnuYGyMFTPMgi1g
uAjnsQeytxz1l0R92BhrrLxWXymvyGHZJQVCFODZKV8thfBvaG9sloOr4O7lRILNkFs8BWT4feY2
BhnLl2LUExZQt3vckLY8T9k/UY5hRAP1lXSvTVefU2sIG+RG4nTkEJDCDFupQhpk9MjOux+M44JM
kATK20GCjHcXxyrnyMqnU699Ha1gfcDaS5F6is8a8QPXR2l1BC9NyqBffXjNTWV1n7/uvfsMjVi3
2ny9oDqtZ1GRxqhXDAbNFAoUDs89IQlksH5HgZiXpdLawRduiWc1/N7ljozrfOIffCFGp0Lpmwu/
1G+0+QevNH9N21BOefhkM9aiFZ33p1myLNv92pYY3UbILAYvO4U4jU2iIWYN2/PI5u4mhVKSVsHi
ym5f10vbwFPYXr65hhFxColqh3zT4NF4RkJl9d2Q6ecD64jFH8U93YPJCUs73B3QV8BYpzMLGlVC
5pQCyF7EC13DpJiva8UbFjS6NnLnh+D1rezyJ9ykOZ+YmNj6KSG4PpGBeV4JvXqepgvXPIBvJAQ9
R/8gjTuv0ZTX9IYeNQ7npvK/jUc3t63GNBTdk2opAlc6vcbCk8dskrKI2VKEmLGyqE1osDhAVYWs
ZgcQOdnYB6oLzTDaglLvMgWuxGGpYIdTsBU05Hwofp+Uv87J03D24SAItd9WlThUZ5ta5QruEqOe
3T2mTai5vDXmYG+WROKIL/buaF89AqIr7+D/4eRTA9ILhOO/G5X3eBI/gIXRDS/MBdxa9WErA470
rX/VrkVXBhfU5ZT33EGBudFW2cKx3Exx8zdqQdfR13Q6emDrjzh5Gm1wT3ITXL78klQqavAkYRrT
ubSL3+GFfvuG1U4R4F5FC0Yo1gzrmzbCoW/RLjRgbaCimq6BEUijhBhVDswwx7IdqJtfevCQWlJF
z6Yi9cGFmQQUasUWKKYe5oL9INJIBbFSv2EYSu7tYAS3nf6JUM44aQp3UYxaJtbgQElynsryGcJv
aAAQh+dNNoHITgleqL9cJoxq0p4Re/Tvoy5gOh6zTpI9nJtQvZR55Yja+TmfaIb8puwsv5FQmPo9
fIKl7om5wiUeJWt3/WWbWYhCqpla49cVQ+s5/229dl5QG5Pzi2qsBZz95hN73PYfOcoQwwIA/i8Z
B7wMHO+U5FG1mLU6Cn8WFWGcfCfqx/i+gmicidYKaSjcZvZmjNiY3Nhb4C13RqPWCslm7sa8OlKe
lxOpXwhVSWuEhsx+gA+8oc7+HsgyAS75ZBcA8D1JoJqhqhT4+nEivHAtg455rrjsDP0+MQqErxqR
GiqnLuL5vJ4elD2emYt5yhgWmoUjmXu/TMDmVp/CmgiiU/6OTYWZXk3Uk1QOk/VnMqCsL9ONtEY9
D6xoRdrj1ivs7OsVX7JNq39NAtwWnLfsCWMyLLGxb+tdb4hQf8I7BfwrE31gIpT0EzP0Wv4JoSVP
tJlYmblUZzAroBNnXOCMDiMwPiLg6/gYmcxuy4N7dsJNmOuxiwZGRfOG4wy9x7xws9z8gQux2ZCK
nC9FaYAY8pTLfx017zbIJ7u7bEk9jRxGuWJuXxKDmAREQ/O+xFjMowQm+0jKQM5U92yN3otKldDU
Rl3X8+XL5Zsuxk26XS2ngY75+jrtaJI/brAUu2+HWsYfa94xF5krzOQ2eQYcGKTRvsdjr9h5xk04
vVbSdap16zIJGaiwEBxmAJ+eKdiRiUP2PnAuKlu6o7Du/Ra/zHMR15X3d3ygo4y2wkL8V1CphQ2M
17sx3OKedvJEIxoiDyFD60KWr5tbheAQJlFX0z/Wn4oBR8zk2C2baZEmFA9ZZT7ZSS+HLjQvqXYN
1OYz9Vx2uwx5z4Zankbe4F5VsJuKynvy7x2BPzKbhGRYhIN/M87N+78iIAoR7dBtswiwDBRaHrVn
s4Rwtj97JNkcVIqolTTJ7YkZwgI3d3fAgUgh63Eo1VefK9fP/U28cUHFnNdMczemXPEUxvLrkgYR
VYrFhcgTaRUrO4VJetDGDMafTqdSrkRTSzZ5VbXJNBE8mUTdiHB7L+BRoGYHV5mQJWjQA+I/4Yj2
/sEhrfA9wQaAj7MxTNCogufEh6oQCY4mzyYmR4UK5MJ4DXF3QYL2IF5eqT6czn+wBW7vSqi6JTjP
AmQ+JSZif2FOuDK+WrkwPFzvVSpuTUFNq0aOoU/Axy6QVqBX/zxtZhSzfNfexFLzqqkTula3cX4U
OuhPJ25okqyI1xpZNZbNN4INIzX27BOQkYqwQLmLdae33c1yDZNFz4Idhi+AX8Vq9Fm9IfaWAu7P
R5/BxdNMe9OoWxLJKz3Uo3TFSOqiDK+1YFe/OK+caZTpRiRuRNYGUHIAyi0wvM391KN2WsGcBsDK
bDu+BjKDIfDG9Xz0507TNWM/2IJeveJFYec2EI4DfDbFnZ8AUvBrfcROuuRsnW5F8oqlHF/Mb66c
FqcR61THSTiFJCwGslY7uwPp8s0H5CmoJEebDRnR5PGe+Z5qIooqmFi3b3eqlAj3ScZ1opkRsjhA
liHNRAeigOww92qsxFruthJSizl+BvLQKaWEu0Y/7BkqR2H6WfZ2U+CCgDzMfe2Cv8PvTIprXgL+
Ezb8urGMAeVOZKfAFk/HAgtL10FEuWr8e+v/Oj3rC7gkxEcs2U3JcU/0piBNLXLFs21jb8OcdNHO
Zl1+HMbzKRdCb/VAfTKEPpEJq63f8n+A5kTVt2gWY97PpbeoeDDfIzmk0jn1I+tLeVaNcqJYiRL6
v9/5fy66AaR8iOhqlnJkQMMeAOeYBUxoED+R3C4+XmquECcJbpmMEqKCR4Wzvy1Ua57+kTDbTX91
dFNI+iZUOMN48PvOS3VhUzTGYP2gENlTmJeje+hmLGdMQdxPzBMRKiJrsRZPtwvGL4VpXfBrPqSj
YC6nhJQj5vO6YshLDV/9F4gxAVkhVvH9HV6L/P2ofqx92p7WA6eWXJJlwAu2LiYOpkn2SxgFlSb4
ODiZ2uXC7XZBHrjABXcjimXI3XZYSHpUUNybDH5pxmB2/jmLB820PTrkPyXStlZBtNvrcbi5FReQ
udbJPQpT0CoIQCpgbl+jFJSc3Urm7N03W6ocP90H3x/dYh/EZt7UY6LXmErgFItcm9asmhfUafcQ
pNjYtP/L+ULdnm86UWNQEel5SrzjOn8BuI3Baoz3mX1iCWLUrN/iEecbOihclxmBQuAaeARPIO6Q
l/zXk4uckhnV8mWPEmeFbFtbxJ/w1bEpYNWhn28zB3s3nU0C8QEJ8pP0QGp68BVeitZzSwMa87+F
1nkRoxqhnnJnC3vo+BW6HkN9ZrczinoXlMRyo72B5M22BbM2Yrogn23zmLsdZzORumvUaniCC6TB
FMwZ1Q6yNqBS9plS015S+XuAfJnoUa8Tcd9vWvJWnfGQd1fYlH/7Fv3JFwlbZ5IVBZ3rrSMyInu3
zVXZDNfPqZipnKCB7mcvH0Mnc96LTRevMuVeMxqhi08IAWmMqaCkM8VuGiBWqMde4m0bAOLE8Q35
vipLa4BUX1Q7HgpRXO8PYCVbco+naolj/8twXKnxWL35VjPnrPpMs9hU+HbLZiPAC6OyVfX+6C+p
sd2oGZoRHvw0STOdEc6EdemblrRQWu57YJtlx6zxamNDFgeALD/9O070dyeEkoeo6/R6QXGxutH+
YQe63OT94Z1eYuJ/s/07ZS8FQLUC02drAytueGL5iukziFQSx6f9nTQ4cvu+r5aZajpSvYyC7hYK
khyQfGLEV2JBrYTDl2RRR+/0QYD+hdLou5Z0MuXZwUMh2f1wIHHARvz1gamcGInXBoKkp8ASElph
CTOsJ8+JKN3XotTSRXxTcZgYCbY41Lpcx1B6GDDlNMuDF9e2qNpLpY8QNAFY34J/yxHC+7BhGTME
/ioOZK+sz+ahZJny/jHXv1lQS4wiHGM3N9AM/TTH0GLuwbi0Gu07p21FWlWu/yAwgnGLS1NPwnfg
+VpLuEiB6kLEyDXZCC0Vfp63c12RnPD5MJrjYvX1fCrbZVc1bvLjZtXBxe3S6g/tl7ftgGGVvBaZ
756LVoXDChm3BR4jYf1YRrkrKE7qbV6vOr8Nf2ZrAQPdFNLdSTtIqA5C/CUzHzzXmFtDxhMhJsJj
io/8uEQQu9t7uRY2sdv9SVNVFKwZPZHI9GRTDIsukP9LOW0a1icd1G/ma6F56wdK0Z1SEBajCdDJ
e+ck81P7z4QR7QvAW9gH3DQ+oca2p2H+uYGxwFT7awXE2MK5n/F0c26br++m9rZ7r9/dU11LUSx3
rXwciNhTdF9ZYeyHRWainBcgqYcwLHFgaMQaGpEpa1w51XroiI7ND5vaYy3hJTjZxjhtOtnDexZs
qDSRaHpgYke07tBM7u3DUi+PGNk7dY5fRnlxKUVMtLNVlp+fVHbWiZqh5zr9MjXqMWSrh6mMVMX8
bGpMRsRwjJg8okIb1xA5TG7KF1re4LyGJLtBq9rtgAjuK6bcO6SJEA/zHS7lX6tqx30Ww09tT7Kb
MNQ43G0TtkykCqj8DcWSYBGbGiuvHRBl8Zix/LsZt1lv1Ln9DNoOohq5KoiP2xDr2NL5h9vzY7HR
Vf6xTl37+GgYW7EkFQjmyGd9NYP5dlm8kZNf7L/9VU7VOncHqjUf7KXLCa9O2fP1qgITPB+11/wP
VfcPgOYuWxgmQTGX8ara7Dd/77FQgJFoI27ssl8zV/z8LPKYB+6oE7EwteuubtmSN0JgZPaJ4lH1
yNAavVZvys08nuEqLimfjM5ap8ZdVYS9KECZaXCKeQFh72rQhWkUIxg7a46VBF4V3hT7QUHOBx6u
NKPqeMQjKDHpLxjrOmdLxlcaXWgfSuV/61Sra8Xho/EvHlruDNx8RBGqcYXI05y0RRTw4w6BugkK
nnw/nQBiZSyOCuxYm5ZpDKabYOjwPXsR+aRezrCfl1ZKhd5LMh7Y+vhW4HuzYD5QxO4u0OvaGBj1
Tatl+YE8/wD7mA0EGYvi5moZi4/I1Yg81Cq33okuVL15yFN/MYTld/4T539yN4yw1g3E9uLMFssW
MkzJO+s/g2UOYSC0zMGAOiqDjMEXPl4F/7t6hdxZ9M0vwKsQ+N6A3Z9ug3qr/pVX2ITIb86Orb3Q
2GhShn0KCkj/5qpDX1gC8ahwzd0wC4ki6Tu3m0D5S5COFs/rgubccHQvsofHTftilscUZ5MwXYgm
E5R7X944qltSqek5IwUG8E01Ar1Rkt19SIylcPI6nN68O2eeFk/69aY2To9TYNt28j+W/rozDou7
SbQR/Qql9klugyQWawHQ9oq46EPRZrCTkWmW+6ljsKhvQ/vDy82LEyKH51AKJSLEKpFex/5Rdf1r
ppFC14F4DAGJd4hi049TteEMyKXGWy1aAKp9Rxqm8vEiBk+hO746RLPy3/oLTdWAHilRhmnHiVxh
TRKaSxeHgRpw6OvuQY7sdla5waxIf797uVp812Op+Uki5HdVe5lQIPPRcb3/+rJ4GsMHC+GdXYxT
IcQ0YLbnz97lyE+yKe9RhU5uM4jfyLnxiVbUQamLS8VR/9g0VDCYCmniG+E6Uc0XpxhLv8+YW4/3
FZds3RVzTDIeJUiZFOq7QWmMrE/6v3Kl5uasNvPuLwhPMgG9gtCbqgX9alD2P9Q/ET5ICBnEE2UY
exFd6ENlg7fN9dpD0Y8foFLfHzKB/XvuR6qGYKrSunR4G9PK1uirjS+Hl/6I6qAdzYf6WhCIp3oD
qIPAqWwqfdIZT+6euqbr39TKnU6+D6O0zcmn5D2bTECsdW7MzVxkZAgg0ICYnRFxGHzEzduVWb6P
ks6bf9R5RqndsuFETUcctfjaSGIuDB6rTtoO3oadm+epmDBUJ3MoxgyiqS/QWzbhxeGRBTeXYf1U
5tILi8KiytcrXUjwNMS5i6Ccc6Y0q61lRErqw2yDd2zTBIgWSKVEJX9WXtU54G5dKTzGp7MDQV2I
wNUVcEfh3uUYNUDeHWt83v59mdjPnS1ukxQdKvS3bLcRUv82J0B+spLNv3xHyiNPZf+U3du0u7ro
t1LNjRfsNR7hHWFv1L775yBb5KXWEk8NXvtX+L1a7pViS7e1Z+HyS0I4QiQoW2PsbL8xFeSX83mP
n0gvPPU51qPGwSesm0iPGTvxQFUYqGy4U6VrVWZLqGzk3Rbp25SlelX0I/7m3/JVk5fzfTzMpviM
OUHovoIFKI+jueotUFB73XBQ+aWdQId5kDBpVGJ5z350tVemyrR0tidGSxvzHpwS5A9Zwpt1l7x/
CF5leBhMKamFw7lMw3VE7T2lvRFoT8tT5Aeh2gzDocgQPVrLs9diBAnhIAv5kgbnRktWubFLCS+6
26O8YS0CSh5VxKWi5vc4EBYoGWrZxFmpDj95xny8yK+jp3jDliqpdPK/7cCu4z0Y4i9aBoxObKVY
Nh07zSlNnfpMzxOxfSdBd6bxyAUuHiOY9RpxNjmLBbJm66c+cBKbpzlKwxCi1DGRSPendoxDgERa
+PquaQ+0uqhQ1ybvcBzd8ZMUve2UIp5H3u2BbD9XpvqulzeAuLNM9ovTmtlsYsfvJg190fwc22WB
n/jmD2yFVZ/gf2jQREr0Ry+W85QVZ+wTeYcDloRU6BoEALv55cPQjgjxKeBDlwDHq9WqgigOthb0
0AquMA/AdsWKlw61DS5BJvNTKXphA9CAct2nefMZ351scFqVyMvRwXmkRSKQls7mt+L3RrRMNdl4
xbttlPAQfiH/Lwm/LqQzh9kIgYRN8ywzh3+4VkseU3T/KQIVQODnXBeDkERfA/QIsakYRnhIIo8Q
N5njgZqwtXT1OZX1pOrD685A4XYV22DWRLjQJGJnwyeDW+PeTHyfge2ePDB0xloFWwC1HRqGupIt
O5+/Xl3Q7FkAZ+PdeVH2+p00FHIb/hiNxlolJP91T8rrU5XSk3vXdyhpn2winW194vfkZaKXMd4A
eE3S1xfrVbuQ30Yja4cWpHWFNUqdvmtAna/C5uaU1OCVGs4ihecUHuV9OtbQuW180Wl9sSe5whuV
j/w/9XsNKq+3BDWrya9/ltEDunuiyzVXlouR6IdRHmG5Q5IPJ8lRGtD+XmCzeNX+wK71d6BDBj28
ZkhrMVhUYmmSxpXLeGgu4mGrtpV+D0PlNN97L7GuO2lEblQDkrJKICeBP3HmpZ48JFh4pqAFmI1D
gBl+zEy9QZ+ZjnT79L8RIUiNhP1yZIHKocoBfUSjKz/54inDTKRrGlj19YYc+4zLXciv2lYRUPYd
DmDgAkyPn5l7yiPLBGn0WjVWuykBTJXE6K1vVhAXRuSmFIFbW4pO54U7mwz7oIIPsdN3tZPw0Kc3
4apmzygZ1vikfzaJwWP2JCKDnxMpmP/j2ebQYnP8kKzCQJu/g75nqNc0D9OqAhVyzIX6pNnlEpvJ
DQ9M0JiS9775Mz2MkIThWmhXdv/Xu5MLud4QiFrmVKMR11dc/438hhQy1UVqOuBTuXMYCVfcdG9m
YXRxaySwhbX83kluzm/Y2SVsH3MpzdxSESF83aTZ1UchF5ocDUo3b0K4zH7n2fZqood5Ujt+0qqh
eA0r1RCiigKkzhLfcbSTRWhP5dttI3u2w/svDYU8gbwzmDZehep1jrz6eaJmW+hM8us0cDNcupnA
oz5fvAFZGh36UOvloLiGO+KrFROofbXceUTD37Yq8zcsX9sCeNI//BmECO/0YA4W5Hmzx84OyJcK
pN788O0XKdMGdowUrRIMHtmBP/eOxTdJA8/L/4jupl/7tP+VWIoq7LDDT6L1qYcpPUoxJy01aX4H
4wVkBX5nYye5jFtCpIkPa8+9Vs+nTXfUQzO81DCeOknQdtxY8iOLMUYeUODqkFBIqLWuJESGQGzU
EQZIja40D/GrH4sxAFX8JYjb+Sk1YxYEJKsgrPTSSg+wtRTp4LJ95YaoGEoAga5Twov+lZKRWw5G
k4dxAaydt71CX0O4mHChsEyOJFZWRBg+a0aKbxJK+Jyx8XUWQeJPbSRVNFJChxjaCbV2DAVvQvl7
hg7M3N1+QwVc5VsLtmXl5MkzXwDHshxeQkq0qsYg7QKD0FSCpYPd7SVqitFbNIBzIlz/ciPty4sk
NDAtuwvC82RSRMS5UGoWGhn5mVkNrYCVRDdX4+Wk/DluMBGNwWLAw8NFbPHn7tZ509GitREEa6mM
gF6dpsshxA/hUxK+pOVBkPUzO4r9fKEl5apGZO9uU/0RlXqQwGJ0uYIl1Ofcs6lxyfnrlTrWxwmI
PYIuGAr54ViLe1lCXZcISZuRdnTj+K6cRuLdn9r2OL8NiNkGIYaj4mBpvgjBio1cyunTSNSdkmvj
KEiiCSnZ6qT6Z1TJecwDHsMTdZK2dnU+82XJNOMaiTvtxZ1MpMyjDK9+BStH75R9jU0rdEdvMsc7
hFyd7w/KDmWHhMjlIXNdtBguphDBnPO6djSK5fnkV+HwqR4dE1sXm3avPbJyFz3uvi+SPLzQLwIu
98zedBSOxk3Thyc3xyZA8sta9q8W8zIaYPxOx2CR4W3PUjOiKN053I3f2FnO6ghKOchUrZ4ZSZAk
97hpHXWpVjVkx3LMkL8FO+ZW/2xEHO86HQi7S1V3wYxpkESJPIFEb5UrjUjWCU2S92/PZU9saLVp
/JeOxeXTW8MHe1R8tHfEn31mBEg7JKRBUeX4d9+MrF7s+ZnLya66CVpfY+QCOIDhW9IMQIa4AOiQ
y9cD3mEkMbxxUwcVgh+mVToXHGiaggCC7nblZwBACEqHUEDthiprtqmYX32f2iBTDxix76KtabTs
9PSbHQMzEsIUjSXj8LLGYGCq07EWsW+IAh2jFQ5vNyqxpssPgUvBjU7w0FA8khIu0hAjjlzEcckA
59+bvaPD2xJfI8/7ScCuGnAG9ZM9Gvfq8oPIJeL//Sf3/GdPlr515xGY9mwvita9CPDHKOZwJ7DM
dxvSqsT4IFLT8m9NxnDmdbE5iVYgviCsyVaSS7kQrZPQtxZ42Ng55b43EZab5tCuVQz8Zva2tuEs
U1sPQdkIZTT1IJgX7Aaz9aFyMrqLbTgNShV529EtWdSdyKGq+kDNGEltLTlsdWWY1WKUZeMbfibx
SF0F2QKPxDiV0H8t/DKBa20tUhPFwz5tyEl0o/mW6LvNaZrIUwoMM4FIVV+0wiCQ1KdjVT0PWTxW
aurvVOpKyh7lD2pQ24D1gwHaYGYL3NcUJz7Ye4+ZCyofWeSYFtvK3SAMOitexNz4AqTri6IRKlAI
SNEp2mb5iRW7S0HLdXT74rg7k4I02M1PBaEv/gIUvwFea8MwcXza59LUrK/DqDPZRMutDis4eG/7
7oIqe3YE9psNJyRmZujroUY1g8sPwsBlCm/e4CUGUZK1m7194n/1TmyevNUuF5k0TQZojHsWQo4/
5PGXnwOZIGN1Kx08ndCTM9WY3xMlPUOPWaKtldECacOskk2FuOXJDcvKK95pulUNaUotn2dz2xJe
bTHywXYbp8+uvziMsj9H1NQE5qwdbikE+2GumNpOyWf60hG9iD3nQEPmjQTSpE1xn/dvcIOKYjPI
B9ZAfRMQTZ1rD/o8aqH7HfVj3s0t8TO8FVOqDUtdo+kVdSCebhf6cfjqi8E93Ep7YcoI5u+e+1mU
TTTKmefp0QWjk+5fAWCKBIndmtDziS8i4y8gZmuog/nkDzTwFBUlQSqhs0peZ0uh7G6cH8u2yQvM
NAh7t93lxSmduW0T3c8zP0t9IA1pvUJKp1kG/UmZEhfbQiIadp71Pmw02Dy5Dk5lQEMd9X98lReS
LRO7sgyuX3ZlRWGCP8hcYfziN8h9WvVxIqwOMx8g7TKtW8rGMOXJ0ZOhpRoFUmfmZPpzAeAV3l4G
4dm3gwlAaKuy52rAibCIEy6cXJ2xtWI86fzjhtmREvhuyoW1cuBJZWfv4io3ll64XAFozYvPxBmE
PRPzDNOkjXgJ2y1jBBPU7Nuc+29di9dU1QyuBpDgpyIo3yjaUpexzL4jFOR5wBrxVsdqPiu4j6xX
DrAbLsK2St28QiS/prvNTPWt7+aL4xAEvoqo960A6Eeqgkb5HMB2HeMrHOHyt/3onuZPbTmFL6GT
Kbx4Jab8cs3Td9cUFMkPEeS0hzIVTFNIGyDI1MYVatU4J5zQEjzCyXp04LNPJZRdKBzXH9LALKyo
3ES3ueEzGFMq9I/yVc+Xj8WWlKTiYK4qntYLpbqu3i+Hcb0rZHIfQLHyRbhfqXy6DC9xqBMjSLbe
ywT8RLPu/WYOBl6wnbkok6u/oGq5EX582Sw4uhI8ufP4UKujojlK7v3VOE/n8/uvtMdqJL1fhBWb
9zQLm6ilYVteUI6aaW9SDFB3n8VHGVvhKEW4KuZ2Xkp3O+xknvhYUClCA3sKngX3/qQzuSRDFm2/
Rfm5sgzurKYmj562GOaYkCXMe+/x3zKHvZeJgB/GJWGojBxmI6FjcdBqerbS7YzCKkrxDB83b4/r
0BgIRUzCmX7oUXsg/JL/qQMZaH/BbgCqYJsVV6oDGwHsUHlf+9xNzH//JC4ZUPA9P8QL+MjUOm+U
nAmA0AuPxJgegTd1YAfR72ETFgv07J12i3lAdpr6+taKbQ778GmR/XKbilth8gpTAm04GlswN7uF
3FUoT5+igW+t6SBnyi6k3gLHdQZnvFP/zuU4mA5xqFw1lVaCcbsq7Wp0YpLEyQ6t85j5mGtzsXnp
gqAyxkB0+Ueq4+3/aFsjZZlZMyDHECyg55KUh/S9dCLbGWFHYvmdnkVO7wimWuU8W90lKRLaZREF
IigG7w/4dzIu7L7vqDTMudcZEC9Ci+Tm3UnnfEcdMm1qq9hwAwWedrT2D3LxLi/o+AtpuGCFjQB2
2OFEC3r5SnnzpQlEqjBRGYfKFE41khibyJx90BjhhUrQ+LgOAx6BPX5tUisHp/dFz3oSr+RJ+eZv
DHmQaH4yDf+w22tK+jNKEasJpteZ7yo3gLBaVZ0k4TKAcXTu62tm9S7J6oT1mW1F1nqXtXJlelAN
9aGraTBpSbmFuOCOju7uKrMmeInBhs56m5X8IxUPAAtWouPInB+gDDmvA4bTjkbLI+HDoHxIgnq6
6P/fgnmvz7QQ6W1E/42XcKSQ8bn13fuxj5Gd/Lpzsoq+9vK4qn6QzO/L3xz7fl7eJiu2VOnTfrqb
CsjxSz94/AxJKtFcQKaJyVNCUNi+wUJpbI74FpB5bn9LSOcZDGfswG0z6WLvoxUVb35pUfMwli2o
t8Ga97BeYQbzauf2zX/95Jbfm3uQ8xr/MidzTJjaTLuMqZCpNSGoT+52p5pPwSpnwjU0fz/11tBO
aD9b3RzdEi65OX1x1EIddmjb9HH3hF/c2yBbp18wAi0cFY3+3Kp1doTYih/AaLK4oo+3R98SdHkB
jhGXYfIeLt0vgTrVDx2cmm95z+WPkk04//8ZudrhX2Fknb9vCyow4ZFw7f9bvTmzReRc8lrVKbAQ
yUtIWMa68ZZF4QfFdSx9C755XeNYMfuKTWuudQ9C6ZbTYc6Twgufgm6N43iv+913kdSqEhUgLmjT
svjeOOauRaZ1RGc7mQfbv4N7o1MeGW83jPCuMOZZvDjLlKGu98/mO61TLkVZi9DhYkYj6jBncSVK
mNAChnnoP+Vrfo6WseffJB3gBGlKDh7TDNdM/VdZ0xNXOqKR+5csOP2zpT60Tu7EawYguDpiWJkf
H/VQQuhkmr6vw7uPBuF5qyzIBuYc1gEQQEis+IlxZk3TEkrEnynIzISaZYq9losrx2VRmUFko94g
QbPujfC7n1uTFqCrme7UIvmTOh9WY+/JRtdLoElTs5c9yERTPCvSGNCuGVHe6T65bCv6wU4q67Rv
CvY2hSILhbJInFH7oYRb9yLb/KXeruRC681biHcLZKb++huNpMx7ROTVzsNypQAP/y7luo2CLx1Q
N45CFRlAXrMj3HT1wNp3MKBW377pVPFxiXLi3Ts53Zakehk2Xo6TYf0usLYd9ZZZCKcZjnkpcgAz
5gm0jIkXcmgehCnnx1bKgB7KgG5xTREpbwN9tsDPVPU3uLrF21zdSDrN4a80XOGzr/QqzQ6hl9DN
83hELPwo8EnPqW9VmwmeFj+0e6g9H7GGD17p95RuaeYRhRiHPreuWvY1tDqvuv7IM/zdOIkgjjY1
qvhRrUEA5E0NSNN5+pg3KXVdqFrb+hqfZo/EpgQA8p9zmpSVSQVWIn7GXiAwI26r+vqz35LsTKPc
8gr8nIwWrgvb1xFaNZ2H6NcGS/Ogmx41SwW6/1wcfiZPOFQNWKmuk/Y4PwXNr1d03akm/F9nIbus
WdSRB0x3nAQ479JH0vF+uDkYIXONgln5kZ3/Jv0vD6T2/ErUkaNzlNdd75dRElzc8b0jVnWqDvmO
WsIPgPcglE5CORdPLfEv/Pq22BKy9Uj/nYNmW2MXQSjjuPkj32RTesSnvEiTLmcSspKDf26SnGGY
PhUq64c0SaGMzVeoEelgQvdw1zmMwM2Af7ZAIUOAnhXHJKpACVxIDF7w8ESrj+FiYS8ILZ6AQTwl
r5dBaj0/OQQCZrBW4/gWo6KMa6Kmz51hY923zhGXLsVW2d+pKCVTrVin8HJv10VagrtmRHsXBbTW
yIoE6iGc3J9s+hXY7Mps/842eUghNBzOHByR74vpDZ2VrB63MJa1hbWlvOUelgHQWHkXw6nON+Fs
wXPdqoGPK/88VlYBmqVVWddEOqiSsKe96eN8NRZgPwRlMTE7dZSAmYJtp0pGZzKPeZOQuMrdPQOi
c2GBhFawM/Y7zJATvOyBaEMmxqGiytlKjg012MDsSruA5XS61owmUXbeLNo47V+YiicOQKZ7Qa66
S1KvEhg6IiMsfcDbhSm/fismXpDlM99IPGQM/gCezqLFE4gUUhyxYSajCQ0dB51eK0kqIvAz76kw
JYNCOoJ9YEd372zeg5egJsgTs1uLnbB7lFVUQWoeAE85cLb1oJM4ti/3w09+rf3+9+jf3lgWZ42C
eYt3oCHZpEaeyIbkiO6gly9neAdKuENhO1knNmxMUbAeiLCduzBAmD6y92MW59c/U/TTzsW9RfZm
8+AxI8fSa1UqPuSLBZ6Rwb5QELIqViHEH7HjhVAAAi+JlZeCW69+kWQNTZQe2zX2TztlXe6KWic+
GE6IYdEVEfAq+/msLquzi3X854EP1kr/ZlHFK3vDg0Mt6/MMRRQ8Qh3xjGkwV3x4gBd/A/XMRVhH
T45lSeplXKV9TOEpHOpruDWzj7eCilZ/m03kfu8I1P46B8yITCyl3rr5ov9hx+oq/kZZuJJO7MFI
kLPm3WNMK2a/9bQl4h4rumLK5KH1D1FiZ/5uw7bA8qHZYGP1fF42PGpW98+fvdJnnaKWWFSHehUQ
X3xHD8HzF6HzulhDZQDaDU2GZ6XQgiXqs+ODHkTMpqiFOoZbm8Gh5Se6JJHSYN1YPDhkb9A2oQdf
zN7vQ6ix8VftSlD/kviTAFIazzmJ3ohP1tXngUswYKsMLFKMj5ubHQd0PjszcyZe2Ho/gVu12i3O
jT9pKeesk8GaHqNraYUtNl0SrP1/MT+fNajBs+4mafm+pynjLrb3PETVtBeZE8GxFdL1j5wk+yAy
AV5iIcR/Tt5+98Gfv16tbj8k4XJgkA+yv4o0LiJZdDINOYy9HEd8PFntJs8yZDEHKj69A06zMFHo
fY4B82GYPm/ZvislkoTG5BvkjF+e0krFlkiE8x7vl0CFRf9yVrrqUv+rPdWJlvi/w8h2YvfIj1ts
T5BRtIC+hkEPudjpoPTwHlVuTtvuTj2aeAvJC0lgKOxyvjsdJhGdf1NpZiCXx3HemkgEvRSY2Tzg
XuWypgg0l3BmhRw7ohJc+qcoAUmw6PvUpQJZ02EhEZjf/bN+L2bBqTmNYIjGG9cy8nvxf76iiUg/
Rrmix3jvRwf4l/tjD86oB3Yp+F22geufFenZTAOWJ3cn4I1IUreMHSCBHLpc7f+iWxpBPEWREawC
ocS7I2Jb2FbSShTYwCc3vyfmT/+NbPxm0VyUhBSR+Jn25mXf0EYD/LnTf2FeLDPiy90JBMI2JoYX
AM+HJhOk2dOlGtpzvzkeNXyTiW+ILYU3ngENkO5FAPc9mDRswCzmMjsJ8T6xbiT5CZFnIXLiHSPj
nt9W6ZteqVsqwZwVygQdUl/AbWUrr/d2vNTPYj27kqaITQ5A1TL3k8LFYQ/PlUGYe3I1naCUXcUf
8yYJVHBf8WnFCg8ccSCJJxH6L2bSnobOnzuvEqhYsTB7S/+vabzvdFZnp99leQUhfw2cSkWXr7Wm
H1xlpod4GNNagHNaPR6r8FfiUTxiemfuCQWZX9Q7SVYKiMNy8T9yAM2fRs0PPkFIBx1UQZ/HbyW1
S2QY3y587OC/oNoU0exDBmjc+50+xs2p62Ixw61aSnJ62C/8+XyfMLkM3KtAjDOzbc19szPXd4Ll
WCw7osgcEpMgmzr0wdW8iOSedRYTU0MFHrnjArJ0hrn2tLAnRBSuHG64O1iLilz5HuHCfmSgBYhQ
lCviHh6I0y5R4TtrxL9F4Dz5uoaoZvSDf/vPGvUtk3R9m9T91vguiJ3P5F2r4IWprcB4KRWoMF4W
Wb+oJ1GxOEyeHlkCDP0iaUKwuxXSnCWCvfajBImWaS7VpXGq8maYuNgW6GnKPoQmT1mQnfpdLhIo
egRUsiW9TcSRrBhdZIy+FzKMD4DKZBQPCUY8Lrg5Sqndgl8eWJReoJ7NSeF93Ymghpv/1Elkw++e
SyF0WrqCv8IMUNsGmE3rkawPgmHidF1oQlpaBv7escG2HGBB79zTAD2W8Z9ImLFams3phIIDwyay
/aFwUYvXng9j4J0wi2hELkRaas4nzi4MR2grBYu3DRKqftAsJN2Bq91pydrbdjbQ//j4ktJgGvbU
od/9q4SAC2gz9MuCb3soAnJ+6qzGpvOUdN8j68Ud4whGxxWLhOFp9OkeoEBlkwh6I8ewF5APkjXq
mjC9/GUk4UEt+3W9tuQuvFw9huTPiUTmd+79FxCBzm7F0bwIWJCfKJiwSZ/7zAPMZmoxeo+6IYvj
59um6twrSp27bhtlosb0C2FzPM4nU/UGMxpw9fo28wXs5yVrnPPc1MynrjFDcX8X66q/mZaga4q4
pqXKNYBTrFvBekxZEEBZvqRM8nAys3BMFQgLzC9vkhsZrfpxaDJCVUY+8B8exVqKIJOJCV4FgU6f
REJv/uFOa10EmkR3ujRRqR4Cxqg2BCUUPCUvjPHDM/8jt/JvgYf/PG79403uD9Kickuvcy/BMMOx
6f68+RAbBcjgSs2lCyHPyoxqJoAYHmOcWO2HYE6kqxH80Gr+9YGa4cGm5aouQoPJSrN8qWWG4GxK
ibFGrY/+mXbg22wNgk0CHikbdGK5aRXa1ICWCKw579F6f6lZVByRo2kxDJ7NVMBAXC+b/eL3d34q
/WaVu1HNpdJu922SOnxwd6SZuZu98SroHbWkSWBwCXSaON1W6xJSUkhdHmXMjc5psB/+SaGN1qTR
8gaMXYLJUfdHd5QWAr/fFWJlUOoCPr0N1jJV2RTZ7TTBuAdbwhqxH7pPPVrYlqdKkW5hIS29qk9J
NNAx89+D2J3+ukORyZEDOiUXa4rKj85c9nJIo141I0O2z7PIOhhKVZcbAzcyF2PB2PaEo1iE00Tt
FZhs03HVlC6J/FwkVqljgsAZlaO4Z44xGwqYQ5ROsMf3EAghk2mWFuZkeSzGBIVyV0KAQIn1AzHz
RwtwuvOmZIbY3fE7UmYoQvk2TVR9k+Tlbg6kGCW5ckfWBQilMZOc4IbidBnlGlSE2RRp4QqJP40X
lZVV/FdUPOioN24HpZHdX6gkJD7JRWgl3S/2kzYzp+GcTVd+L7GwA8Jtbvb7LoMyrJ77poIqGBSx
wJ0DFiDz5rli2+eWbZ7vUZg57hsXieq3v98DD70a3DUD2pF2ryy4/G2t22BnellsWTKip6O8OMHn
qDb/Fb1p0F5VH1Yxaa3jsRzhZ1PVkmu30ql6iG5bDOXx5LvadP9x5BzQRnwCme+K2QwRG4yCeKT3
XYk5d81eP9HWZDR1AtfYgck47IClxYQiTtI7pwkN6kezt8HE3gdzLtuAKN39542TVwt6n8RVOhw0
3EoAkrjoNuqnbT90eot7MKPUt0InxeTjaYnExGBmtKCAH0+LO2PL/TOOZdYoAQbWZ7rP7ymM0sIS
bEf7joULAcZTmPpi3UYuJawTq+XwYHT9NgEZoYjinF1eil2jiG3avFTRcAeEHsJdcjsxM1H+1bMF
AX93wCtqCmQvUVSTi0bYuPPgxJ0VRpr/e1YQWVOT4w692UDhDLK+76baUmqtMgfjOvDwD8gJ4VA6
XY4kKyMPk4xR1TVpuD0kFYqrhxwIapPKcUAHPrFtoKYgIef+82bzIeeGLe1s6d//Uy315aIDbB1r
Yd59ZxpYFrJAjJiB66G/Oxwo8HHENbyfthdZRywAOc3UKjyNG5viPe060caKGnQzGhQaR8d7/bmU
pU47OxrrWMkK3+FJhKRRAvrbc4R/JfhASkbeiDDDI7x0srp2X9nDSL9Qs3esextVakjvTI553rYd
wotgHfPyANE4DS7DFusmxyRXp+W2Sz8iLMpLn6J3YNy+3t0goVicdT3wlLv3DbW8q1NkW3UBXzfx
K4jYIjg9A6aSfU+k+Jrl3KPFR5cwPy8HbMtcqVwKOOrYaEnvCY4F6PwHtQ+rVpUnALB3B5Bk1XHQ
GHlCH7LkDuJlvQgnV9Zjk2g+rpg1WzNO+uXXubpztFGXCSox+a1bhhgfXE2ItLQsUCKQijRL/rSN
CMFT8lRVAiyu5ml2C/J4wP09JLm4MIhUMqMeduDEFcLrM6qPN7W2E0ejCNeM2E8hYhg41cF3j13j
+Ed02DHUrwpwtH5b8mviZW3Do4R8qU0OoQEgTPFfAR2UbKIirRvu/pVGDf5FQavotDqiWrTvZdXd
qworVjICMrHicmLBYiXJt3XMMpc3xH2f/mGAk8VZ8IjLL5c7BCyWfuf9J5cdM/30zojcoiKkdYob
7l0hbO9MlV0av6OXd1u+7/A/cFggtLpVMzInnHlVyRZFya5Tg97Z7pgjxQ9fr0Kemzfq5XLi9fWI
RWFLkKVRxGp/PE6T6bIFFnTJNb/C1hfcV5UL1xzAvO3h+tgGIWqvKGmgyHO/Y1N3b1PO0McGcCIp
ny9SSUEb+blg/mK4YT3SaKg5i01iU5C0Jrz5wCI//wxw+04HH3tCjj2LJlTMyLTbrh+aUkdB2Xp3
w93JBwGMxicVN2gLkYy/9C0q2QeXlUgNg/y0SgSYihuryKsi/wWQZj1RICnCDfDD2gxFExV5eIh2
CAgBM/WKqlwuoEAEAEsu+A58VzHzwZ46ByUd8uEy4bt99n9ojTf5PtUj4IrRWuxCknKAS4FDqPBm
VQnn5oFJbv5IEf3fr6ctWUWyUxvGQpkX4+Id1Rz4CW74rIIEsOi3yjsRThL8+Fcb0qOGjmBZAHcL
IFaHaUIqMWPZ7Zkz3tfzbQvubJrOushEVgmdM9RSlBZAHGyISAiZbV7+JlvT5gt7h7FK/DvF5/up
Bh30wzIrcyGmqZiS4saRjy0jlwztTACjs8a36XFw9FChmsRXIRg6vwcnS0WFsVVDg/eVc9IxraXb
jCoZBTnhKxxIX4/rnZkNbojDm4zcGdCAQ9xnLfqxHp23nyw1aGLzQnpThCoxKmJTfwuT5gxm+3lL
saY5lyU5YLXxK9yJh8hh86DcxUe471vyLjIR7YaMKp9AjAacr6zPAjri/5y5FU3OWmgYUdijW0AK
49f1KvVM6BvpVhspT79WULkbK9xCOrEkTti+JQD4lzQLGUTSigxtBkqszfriKjCV19iO1AjbBs+o
6nmtPzIB9mfKjcyoE96TR0yASzcQhGRVZ+rh+SCgALOkPcpFQemOaTWfj+WqEljrfVm8ImhRJ9zQ
Ce2PLaxKSkdqWcWqqJHnz4pzDXCQyGdN7XKFZ3hCtn8tlQFsWNONwDLSFLfs9v2KRs3lX1q97H7i
XIF2DcgDpTze4UAZKHs4IKhTFKBv8bNy0kcfXm7eTkp/b1Zhg9Lc3MfCKAJaG0mUSp8FDKCOSUfp
YaFtvkFwiZbIazDc51YQWSdp7LQo/N82HHNLIQDFbf3V1rHPkhZ40B3ZvWYmMB2Aec32UC3VwqME
ioa2kOndcyKzjgbMd3ChiYGQ9K6ocmp21ynWe/V2TrrCu0gbKi9A9jRD0ECxseGz3u7nj1cnRx6V
wYG1vYcnbh+eUcnedSIwnuzILMe4cg+yQSGND4xLzA23pV4oHyfJ/8F4TSRFxvf2w9oCs02AdV7C
h+6o0EL9TgLS45L7pYVadupxOK2g57L4YrLVkaUL3jUiO3Xnr0HCJWRsjxaq9cK2YQ77FEmd+3Qv
E+rTAHltpknEw/D27O6PF5eyIgzXLZmvMeVtBxqS93If+iG4IqdOpbuVgALMKHFZ6yCJf9P2FaI0
Cd4BcHltZvEXSEGlFEsM2j88/0U1af82iPRxGgjF5DYD6Pc0W9aPR6ek2Bub9M+74ecDyW5Ukiwh
/YXjJGtMoIyakGwhR7q1/sYuPH4+W3f8iTuYieVIcj2H/sd3Fq8J9KVLOde7rAgxZuJwfUK9fDOd
OPb8IdfPKCg3F/duDSdjRVFb8Xrl5LIUAizgYoVNlZVh5g3OrxEqh6f2yWfrJyOB0WcRdtAcifI2
RX7NdTm3RACv5SS1quhwnTLDUJ4SZ51m1/ylXruqUsgYWAI6qA8ZgkzaMynhz+w4wgJf2PGicE+j
Tx1k721QODFNOOdQERM1+KTdZxkHorNcMXKw7zFXq1JROpp2RlLMXFw9+XjbYHSu8pSfX4kc3SuP
DNBLw6cWJqBxHkgVTb9Ld3+fviXsfmf9a8Zj7HIo2fimm1BRcUBEJ1xk1qd+YBhFMxBaKKteYnBW
7KV4wCoSUoSdhKjJXnQ4YT3G8WaO2T285zCyen7SfnfzZ1fy41YnaUzSsWQnLcIEdH17j404gxlW
bh4iwchRdgjYcqUEqpmD8qgLIsmItWC6yQ0UYxGrsSXyfyFG+7GOAiK58Yvvy18m7frGFnTQA27X
aYXP9nCKhGAJFeO2yQduX+CxaoO1alG9IWwU4u9H2jahv9QH46DgMevFH3/yUM0cc7Iq/EQ0N7pd
BZbIDl7DbrPCcHfVAun1mULpQHQvUhufVKOmjiT1bhfXcpA83y0eIwalISC997NRoGdbF1BblwLC
tJKdCyQ4bKyKG2VHnJrrD7eGE/QOsKvU3PsZH3nX9i3sP4gFmLmTi3nto0FhFd3Of+a3P5u9IXsY
yYLAIP2Q4wqBE0j/CMrK4VmKUevaDWJem2w1rSZXXgn3XNmR3r/RM/7cFBMPsAmPGwEnI2rORrMM
3j/C1NyNdKZ9d0qZw+1zyQxiCPnq9oO6m5NXpBEpQL6pYYW1g3oYhu9k0PQDs73D7bsgqG7URMcM
iinZxkoN47fuGdFnbVa5E4DDuJBSXFO8gtv1yvyQ9PXKV4Bhpn30WQshNOUxS6Re9sbJkhVJo8iv
ktIhdffNYqBRd6pekBut6yumNmyQx0SESaTJubdwjVWyScDooWV0bTFrv53lYYGNr10mulr2iBYh
ISk/fvqqfoJZ0DEBB/ip7YNTcKUpW/vK8MdwvMIYB17Bs6Li8+oyKBjhbA2NTbnzFwuUxRWac31E
8T59h+DWr7/2uRxwCdmxPti1Cxu2fhAqnYAoWcGqZqpfeB/Ek2TS/hCOSZzG20ZWYLCUw29VaNVl
CBDuFPl3UJOeXm134R+5VCtJ2ingmlElQVqi8Ph0AhgXoaDtK6u8nPde3lJUj+BVvKJjEU5oL1kL
Uxws6hemwJHcBW+BwDAh0dZB4mZReR5XUiCXyI0HLzc8q88f2dckiN/bKIL0wExOKRkdbiu3L6ca
cZdGhYEZVpZ31dxdQ1P24PB8Ox2hn3ULKE/l2vwLcp1S5UsT8IBHOM0UKr2sFeiRwqOAx4ysmn+R
3qaIZln/+bfy9odFpyn9Wa/KjpBys3Pwsp8ugalQSoT0fTpwuSBdfLZ2DCRmUk2x0dyEcQBEF4pr
mApamObKpDlat5wJwP6TUcLhw+wkf+ayyZ9VH3O4QaYRZih/bCAXgoO+xsWwt2RuOmd3gfUOw6VS
ipsh+5kZCX38S0XOuascnhgFi8P6hIc4zk1FqYKPBTM3g5od+j+yHM69VGKFuH+g4kvj7EsiRcPv
663VRTXnGn+mxluB903D4Zf12zZRr4Jh4aFOmWxNWnrCi2WT9N5XYZJktYF2P3Ocksw682dhcfGp
w9gMf2S2l42mnh+R/PQIbZHyfq/54d+TZSiDH4i96NZ22a+f/aZVJgXxCUyHQfQozEgsawbtw4YK
ytvSpGM1RvzjmxFoHBm3xiMJ6/ZlnToGTNOQBaW/6civuIBgAyRpBhHLx3PlE9imulJVkdXB+rmo
3T9Kh5LcH+1DUJVie5SSlfbYwxDQ7BBxLBZJCZcy0gpwiYOjcEL58ti1IwWMNXoknDW0ADAow/2x
T4S8Q1COomLBWQwgbGfMLYva7gvjcxHQf1/pEsR40upigNBpepzGtqpMDjSJQE986km6r9uoqjml
kC7peHODeWHC7VwER0dRnP7D6izDsrFAngleNUUNFPC6BTXY2c2sqA/gieRl5g+beVGA4UonpIk2
zl3JnViGj5asHIWjLcEdeCKTzZdEtsyvzRhLxamB+5vTdUXByrTzrQCXqsTRCGQj9LNrSPbiVZvn
RkSFJgeiGRfy+ReZ94uGkGevINIR7GAij/+eA9gjaVQ+4RSSLwryw6+/NDES4udJ68Qtd0uRfTmS
2wWNsTDIEewOC/1Ydd9sL8On3DgosqW16s2TUPsyXTQn8xZlGtmyOi3D1aTcuT27n4J4iuvgwx3Z
drUwogtlLSnIIAznz4/lJvhNavo3puDIw5tJvD/nontqcOrTB5nynv5DpOCNLLfhCpGq7Dn8ZMJs
QWNruLWxJh4EAvP63OJ1oNwBMA+NRSYwXyCMn7sbmu87XXOsywkabWRrqgUr04ZRn12FMas5Z8/X
8sK68lN1CQF8cA7zNuGsvsNxGPx5+bNA0c5AwC+W05/27pAtDlvD7Zem2uk4UvoA1rhFqqQchzR2
oy9hLnllD1h/uGioDcJG/CC3J6/ub8f9vaUJr4OAwj2U69NiHvh7KYdiJQz/PczZ/tFvQtvZMg3+
FSBaDSlKKM1HyCxzyrxx8HNIl+5cxcOtAGj5YFiN3wvBgfPVcCfHJIhA5IfT/exKsBTI20MXy0dE
fsSTE6rAdvS3inSMPJAvUgW3z57Kua+pM7boFWYoeAaNvXQPfxTjg0/MUXxW+BeGX7xqlkPooFtZ
r1oNFOjKG60qK/uZrS4vaLUbC5/L3EOYedxkY2eNYiLmRRatuPvSbsBOJfZYTw07PEDCUGij6rcF
uLJTwYnHcqhpPZGatD+8Myudjs4EJAsS1aP7WQPtec4YNJdr57V3OoO50paPPUm3XPh33VzD56Tg
P2yvCbx/rNAoYeGo8ZV9di9w7mC/Co4ipMm6Eu/AF9FyIr+roLIEjHH0hWreNPnJn0U1ukiPBtPv
D6Qu10yvyU43O44Iat9Nxr0UurqklO5ZDcVd4GbsTfvX0sMJBRbALWPnv+l4Ur4mrPLBGUBUZiAh
i2Fk+J8Qk84h+6jfBUQcGoSe2DiuOzpHiqXvSxQSmCcR8jdDZTTwLXgawAseQ+tbpZAYBTuUhdQh
FxMom/sefU4d4BtWdc4v3ftTi3Z1hwp/y0j1+/TRrA9dsaNs5LGkSR2Mls5/C6UIYVm26TPy+xlW
IzVmvNphzpEnxR2/8Ay+LjYRAYS35Owg3RFOx1xkgoKMaylzs8Y/kVzO20WNM7/4a1gavUHTVjGT
xWC8oEa6+YBov/TWMpDlpBk7Pnbz2Htn/ueZnwTJrUwXa9sAsnfO2L04t8VyKByb3bpwsVzn9grD
GMW+R+tdY9yrZucuB0Cd4NvO+qT+q1+8FRKZmvMNGBAglbzeFI2Mtwn8/1pohZy/jNPUN6RMp2Fn
glLnH8+v3zLNRHF7kAxY633QlEWQgCiQYsqYKKDsQ2mLaVQMOFqL17/LaorqHU8cYC1iX/quPdNg
A3++RIgKbGnk3xUQ/2cr9T1ACqdr5Dm9obt3yYhxuOfEWm50YYqwXdJhb7ei3sp37dYpkdxaTgCI
MtzgvjAQ3OqanGL8W+DvaS17f77yzc0ZdUL01DtubB6uOcahCbsZjeTEVhdlp3Wy82cvZztO01mb
qjJoWCoCEiTwMMxuVSUF7rpirXtCswRjSkZS3ss25na0EoMSJp4rx8ieK+x0lGqJEdvnrDa5EIjK
pi1DCD/uCXnxi82wSKtTGUomuXn6DISjDeq63DwoDUeVH3IpxTgnBeiOEunhBLo3rxTdlIzSEW4l
XGn7I1G7HfgAFJzjJLEZ/QAeKAc/WzhBkTM0TjNHt32sSY7kxgWcnWktWP6GpQR5p2iw/T+zkqde
TODaYPAU/IxnLwn83wFIWvH86vTcc5dtbc7V63iukxXWtv/F1q+E2sQNR+scZGRzllmN8HYiTe54
qh6sC0UsIT48IpjFhhI6yfDEhYcf8SA4dwPqHJy21AO4qYBQFRJOQm9hp0bnipLIgVD3PYtriOgD
v3x2/QUmvkT7kuK/6fwAq3z9KiwLZuqbgLbLRZp9hlHgeb6eQSve8sLhCdxiXBwak9yaa5uDr+oj
B1ynQAX66yNtUlGAPDaUts8USAyhRlFwKeXOpzutqFFprjs7V3hGShUfmIMJdAJqZz8XASoIagjG
YBzqtssvMKJMHfByK1mL0gDIk75wYXaFxkbZ9czaJdXrtAi5pFZxiza9bLWJsoRzhccCB6EBLlmR
ZVOyd/hkPcF0eJnZTfsqhB6JKOXDQSso2OLG3gQuoV28r8Mv8ngYSB0UnXrT0DuLFaT/Rwkie/h4
112T8qUTbgHr6Qc7MrjxRWStQIfvZlP1g91Ny0n7KAUMShf3oYQHK+VGGdnzOlJjY12HNws7szU6
Ai5FKzQXFN+P7PodYmwIFHptV++hkWNxOvoOWXyS5zqkM450YgNBb4gSryN9fcpnYk0eshsqthGi
4dbUddGJ1TChQMEaUMjLbAY+rHMseV8QFF0rJbsUkQlLVK51ANDspaFfCE7EI/BXhnG0k/5RqW+P
S/Iu3o03xhAA6AAUrhd1EkbWec9DNIFhONI3DMGxdQc+MbdsLqt1Bwt6K403pI2i6H5QcS1gUf8M
nh1CFVmHs82wATxTIqDohXp0KVAt7ofnZmg7YCoAEki0DZdcMXIeEbhI3b8iePvXg2sQKO3Vk9Px
g7xUUb3LV8yqnWkEntj2OZzTWSXoddz6NOVZwWZA3XIGj8u6+x+0dWZyTnlWYe4Eb75VAgHqkOOg
EUiRJmYtY7bocA8C731VEmW1TMjLmMvhQTqHAY6bxUln4EWGvNpixjtmzqqah6nzfZFDSk0UZgk3
mO1/0XiVBcgFG4Yfjt0Y8uiobhwCd+7fkaQWiITe/CUoy2duZ979uAJQDg9JqqS43y8F6GO8Pqqr
LuL3iVKChizpugPJykutR+2eNyiE1fjUlFeLlw3zVJJQGezjq0GQ4LDcPvTwsRHdDa8p49DVrsAJ
21QEmEIlUtX1xWylJcv5mrnegOJH9yRq84aZEAos8q0xwRKKXnWJp86QaQvywBhS4PFMHtP1CPfG
5aEYKa4gaTNySn9mzLLfHfCf1AGlQW6NixJJ1yg1YZR6i4Y3LdPrOPAe57wpD06DQUa8WQW6CUm8
9WcYG6RhivTnqf9Swj+k6xcctM3B9PFcGAiWooy2QHFA/gPjh6C/ASMvhNFpTe90qODGsU9mMpi2
MGmUnQ+RboJHvXwXTDp4yoPdOUUSmL0+CxjaM7xaWW+I4IVMJPVid0+UsHljojXEUAutVl8gmxIh
1WoBlxwStIg/onJOuK+Boj4cqE+jvxM0Q52/Whk7nNYYnhAB4JuNXdM2MENOtCEYo1S0dusHXeRv
lZwLjhZ/S/Tc3btmw7yBLB3s+f0X2qMPel8buigTzFX80NU2iM7/k/fKXk34ao82ej8JDPTXe8fy
Cvsc+oyy6mU9f5AwtKC4vl1M0FVjFxbw4D+GICt4cJ9VtqzOx1JTO6cp/thRTqgx5UQV/5RY8Akn
H8+PaEBV848vdEwlelEx7Z4X61c+dCtuMHa+w/Aft7miepOwWOXgI7Wf3U6UcS6ZblC+x6lNhJv0
yXHC+uiL/20dqokOsjkxpNQxa7l400bDLgAHZtqs4tVqKLGYEOVLTFbBMyVJ2KfSfUE/PtTXBJzE
pYoC+Z2uAt6AloAHUwTwv8nO/LiUwJQHyjfZw7sT7pe2eBUW3OMoCitH3dov3eTh/MnBEHpAA6P4
LbediNuMKnuN7Lini+23Myzk7MQ5v51YvFRo7nFtpt8qmlK/CiUnRmQsXKN4qgNJ+YzhamG2a0v9
OodI7gSWswJlkW3tIYrfgyKIIAurYUf0iXZvCn8y6uxZ3rYC1VV6Pa/vJPlx5qPpuWR/LTRj1d8T
iRXNythHfUQZtkNBilFNcznGVwDhcBMySRKoCVIKuJNgdtJxjpPbWjYzwKIddrZyRb4XJSGFWAbE
XuBhLhwwEWOaX62U4z30yG2JsSsT7kaK64lYKyGIfisLduR/QW7B6ZySxJh/ubh4ylJHw96fikQE
T1aLTsjWzWqbVYUW8l6iK/PRHoOXMZPx8msYkFoEB3y0cSSrM2CYgZGD/e7krjUGcTjSo60cAhwh
bC20AMQZZPPTcfQB1snF0NfhUkBjo8KeQ6ZYWUQ3CoxlFj9ZZduHC3q7mATzQKcKW1dp7Dbe13OK
m0Muf8/czMoSvf5Yii3RKKNRKzW1FsAjDg1oXaQk4rUgQhalNzZAbBVyPpYmklwHafXueOf5I19F
Lc39B/n3gm/Ham7F0Y+iIjVSeM1Zhd+ulL3M0lBHS2luh/0owz30etMp4TSM75ZHad+Y1rCSzT6E
2S83i1iJZvbjUI+xs4XAvtsn9n50QlfQAhOmMLUbT1wYEnYAyMqeq9teLOLHr8NpvED/WXnpcb9J
LOT7dPOUH6ppkjVgQa+r5zdWEqfz5paIqrZaEuGhOGw/5WSlAnMBaJwcIua/4tW2+wcJiFBGVkah
D7R5ruR905V4cS5wK296WPd6vpUjbyrxCX+e+nwrWkRe8dEmCFjB0l5CjglYww4rWGFbx2mkpL5i
bguio7CpX2q7ECElL1KWQjRhb94K0vu+2oAYirhJ2cRZcj7BuBmgjLSqVvsVh6GA53L1+UibdKK3
wjP7f+6NKyDXUM1r66gMBD4JbHWuoVg4jpb6wOEMfbKpb9OTADK32bWPDXOxsk0VxVxWzAgEFJfH
mKnLR+Ds3Wc8yrTADrnW5U81UKs9MX64LyGfLv8el8YcYygGnqizPIKMQ16ja6ZCVLNmAQqwVhKn
ZGeVhvP55uiUbUEcvlr63+EopTmxwEtU6M7766Z3jlaBM+/1HxjbFXefKSmPlgQec2aFBP2izmSh
9YWbZQJ3AuIkOKl0xSfMPgnr9JJkvY3NNd0JKGZr760MCp52m95M6VdulwjuefTlGrIb6tZpg8Dh
JyaBM8A7itLmTCSKgycw1TJkOyekkln7UAdSZYCCSJl4vIMwvNPz5WixW1eseDIXRj/YcVHf23Vx
f5+VlMTFQDK0Aq7ivdFvWPLLSgbZaF8SkTwXl3T01ntxcDd6AKq3zmlqlNACSqiLJdfSvqm/+IsD
9bvSHsfRws/etJ3UF4DH0UH0qJkd9Z7rz7uXMDv6ctJ+oH4Ung10LfelDeNONS7FJf27zM4vB3aT
hYbiXvhOnQ8+4+UUrttJrkiyXss3HimngmUEl3ab1DuQIXIORB/Gy4uIkcUDTjHiGRig8HBvrGW3
jgfVeWAGmt7hEK5dvr2akGpiEnlV2LApeD61Ntx6e3w3rD5np+aK6ucggApzTWTL+JdLtNvT+amT
C+kVOY1Xua16zM+lz8pc03zyIBTUpZummHTZp06NBhp0lyuqASuSZ8yQFjMRHWy7DF/PDykkAh7N
BQA9B99HN633bCixNk2uZ/pxhDlG6dq5hSqwZPDJHHBmM6FQR+DB/TwWHtMgKfJB4pvMwDgTe98l
N9smsVVxN5B+RDzGbaXF3ayjVOmn1kGIVnYrq4Wqz4jaVSq7aJr2Y3rf9TPdKd5STsKdrLCw5Mla
A6Wz/J45pIPPoBIDsSJr5usm7HZ8QRD4OL0hcFjkhuj1UtuwI8rV0E2kneBR/oRJR0ZNUqAx1oky
LKJldvwvvGuUAFQhLRIj/kMFPqpf/q1QfkhEX+dxABZd5eX8ytMpuCi+2pSHq8etq9mcV7pRFhDD
15i4jaK2xl744tXD8ob0hOJXfIcVhogJHioCclRIxtD3585+9OTtsUhDHDuqF+ivfjC7atGwWH5t
1z2dMskZsHv57EdUmminENOddV5haba6KJ4dHolsZUWfP2sAiYRLXc/6+GDdPo94tJiSCUNbOScA
r02bK52bXxYXuQ788c4goMl7GI5kFjrX27xDe2tFSd2i0nDbcpVQa812oJto7fsNZOpezJoTj5p2
PDn58d+RN5l6q8Nm0cFqr6ZOtB/yg2olyw6JlOMnsiBLTlOdOX1uAoPyvTsa/a8gpn4KW6fXqkhm
rD6CTXkzcrj3DTau/inhSZCK6rUNlbK/RHtqogX35P0Qrs3i5ev5OFSJNzJyZmKahw/VGzNIsQ9X
fouMGPWIuRS3nnJWJiwLHZ8KkXmslVsbO5r8tVOU5QJNyovXa48nAMfMpakxQVL0kKwDnVcEgk5C
afu27cCTX3LLs3+dAhFRZ39SpYuAFVhrZubLEG9FVZVEH0CgZMhnpTOYD4pw9L9uS9Amnb4cOpLc
54g4oFveojMoAM/HB5hFDk5FoYrRfTVbdA/S6dO1KTpdM2cU2OarzeOrKftjIqQDFjhWFV5MYcI7
v3biioqxKMefsdObSpQ0/0gbrQALICHYVQPlfEB8UcYHjFHZaIkscZGY0CHgF4CVNCrgR/R4Reyu
BNq8NsdogEBnlfVyGqmRfwCRXB/V650KGoYHMX4FiU/T7SC0GU8JbnPU8GxgqN9q5UcydQzUoCbA
tb987D1xb9Korw8M7LxCs6wL/dzC044bONfjcnmtdJEO8TfeI5/MM7VgJPTyh417UaqXieOpbV0J
gb0cHUCecuRVogNxppHdgd31ul6F6dc3RctvaV1F9zIg6EFObokQoOr0yLyIsfkN0aKixJgTgul4
l48w0jFDu0XU2utg+2V140jj2od8xYgLNIxNrkrTzHZdF0oD2VtpIIUBsz2znGYkDX/LGAZ/wbt5
CXw4uUpYkiBT9xQYc3q3Vi5+W4U0abPN0X1Bbm8rmRU80fEIil5+oZd39Cx/4nlfpd3dvAY9sIww
OPwl7dIKNQ0tvpOKZVa6m7scN/VXrFBDEkTO4iRMFHW2BBewdEfoCZHZckNmthkXWoqXHP4LoquP
WBh1j1CzefFoJt8pgfLW/ReZmi+xnDvKcnHg3f6A9cV60+9YBB0K5I6x5+kYZ+gDhwUhcMeyobpQ
5tpETS7BmcDhJnrd4BG6b/JKz6uOMRkh0djQ9+gLIyYBDB6kB9UpydOIrUqcE1mxYT9uDfhU0SYG
TGhXR0YckBrhvhdi4rxgkl9CSESsBmF67jmaAJ+TvIeFGmrnmLpT4opTHXkhym1a91AaGeDJWfxi
qcGNX2tvGe8gDMqZyVzVGa/RwWZqPVeFcPZ/0/H+2kBZREw21ZlzLPDySokEkYE/3sVq8MVNOEwp
LVg2vMBszpz0zlLAlm5FG7svErtsatPDhZpYkcoqYJ54SsFckFN6wsA+eb0TdnUM8RqqxIIsqe65
Y5tYrlWQcCO8OuSh68IU+MXB6n4vysDItgWSr9GouUVaXm3t5o+A6wT0pp7UIAtIWarOq5pMjcEU
Aso6jJ3Jk5jzWDLL1LjM/BqE7qLkLgEeAdqRGt44EbWfVomGsPoryWMmeweHIxMMXzkdx8TpebDG
+pVCZDpyLKsGz0YJPqRWwv4rCQL5kHgS2fot3Ztq+yXjfDhPq2C8tftD2fl3HSy40H8Cb/0eCOew
wbdRMHjjylIr3Gs9fnrVEZ9fXjYMzQC6S4GzrNkCOccwkfC1f83FUt88OzTUaOh5hUIUjVA3ITFY
la3XfhtC+VSLRO5IlQVdlnKRQGD3aGpa+sMl56fpankgbIRJzgkZgbP5BDgzOLaNEisr/kr6HJHk
dHHE4qARFaxNu/ekMUAeaeAkB4nwLJ1K0zqpjgjYHoye6MT6oakyz0SRML2/CkFfqtacmmeMuOU1
oaWaSTd0snbDKtHedae5/GGtLSoXKvxu7doE3ssu0Xr5gwwkNd9mHQQUTehFFWIi7/dbcNHRqGw+
rXJ83bK+PtmKm27ReK2N/pViBP8/Z+E/p4Ch62Fq13A7qExM4CAC0kJvwpIVntFdQEj9vPLQNsmJ
Oglb2jZYVxd1BDItSM8+jgqK4p455lTucCpWYo9GxkMM5WntN5d7sVe1Xo3HCm++YYBWS5aBVSr1
958RVWVoWTZgYAt7nBtQYRMa5XnHTY7iXwPESGLVBzuyenitQXCZsdTQeDddUP4A9AYuZKZsg1vb
bUGK59hyGGbZQWbjBBCDu+L6h/k+eNm+Fo72yJFlDJAZr2CVGQ8L+zG/YuJBM5a8j65XyDfcMsPi
YROkw9cFvvC9XYaskixJM+bYDlQHnMZ6lHIhCPI2C4AF85L/JouwPNMOoiSeGvMeSC0UbnnmW/Au
aWtoT1Q8V9/JBqhJ+y/ssUH3WKphnXsTxFj06IPakBz5pjlI+MDMqqxNejbRQENwu2aAoJVfoykk
LdiIcUjbhjvkADXR7M6b7yoIFlYdYDKD3NnzWgppUw/bJkEJMyIHiSlufcdsfV1rMcBMczcJ3sWZ
IbrqQXJCQ+ZtgJs0S8vvwFoime9/J9FAjTkEhnZCVRyJCLwzERITUXShX/VigVf0t2TIv5/iLlLV
p2d8Gkc176vMoM2EY8tyr4aquLMgj277Zjn3Wiyxzyc7VYOU1lKxoW74dl/+93wRfmTqqxxUkbEM
wrAO0GmsDtBKWnYKkDSn6dfN19TAx7KbxeRTiqwDRjgZH6j9o+MY9U9Zuy4zmHXrd8QC9POVmzHL
/oEGVgg9rjWaqJ43jHVrXKPNUj8DSm3/7SJI06jqmfQeQxW2+yrGtE+aEhJZR6jZ0tbVzcFw+97I
+j60dzIValKwjpfF24Np6MZfRdvLAKOnwibk5vIRW8eXXj4/rnBZCscJD1KQgvzs/IrE5EbD5u6d
YGtXxL5+W8Ld7f/huReUggtHuC7wvaQrafnRFLIiSlZ8Xm4B+Ya9VX34f/SM8POCu7jwHKOYSbeQ
Tqjm2//mi0R9LpIZ1a+ckw0zJArcWJQQs+1CluviRztWjufVyNwAaN3jurnPrj32BokGiRuUAXjf
wmQZV/Z9U8oc/sPd0XBLV9Cg4yIeY90M9E8s/NbFhBj3k1CoycMZAU4uoIq38iXfm+zPjrPNbAPw
I7k0MbcV1G1uovQ9mN2USUPkJb9LTlL+IhxFTNr+NwAakHw1gTE8Kr2DG8e8bL8vZG7VHsa+xUgY
luLOz4NKMMUuB+pOdeN3QKglA3VXx/ZfQfzc0ILM/l6xnmNU3sepJuir1n2OgorGSD1teE7bTS0d
/TQr94jLZheeOblxl9Xapz5QZB9uguyTeDZXzobrTuubdb8ye2SFtz+BlBPzRwnUc6dEzhW35+52
CRrc2ZcD5TjwBl7mftHcxMKLPCLK88uV/FgrkGuvxuIz8HEe0Yx65OREWm156aJ4K5EJwz9sXZR7
UEkOPYhywz9BBqTRDfSYild8xUZKnz3vQy4eLgM+ahd2dgEVWbiFG4e710LM5dm8e+D24BLOcKTW
AIobN8k0qaddyZQv9TdLCN+zRaf5aetzpvpaggGLQ2DOG7QvAw4tYdXm2KDO6Q4pCBBPZ0Uxuzid
EbFgNWRrhmDIU3xjLCjr3elp6kwBGtN5vcghhvTQdWDC3tZdobgC4yL+Mds+q0jvadmfIgd9AUBt
1PEq5km1iUHsSPOnECzVKH9QRVaIAlD24Y95U+WIuyusi9baUbVVNLeRMNckMl4hSm4lMvksuhpy
CR018t337O9rvUf7tD+jxFEHzJ0+UkgK30xQ5zoiPXYEjBP7wogShJeZgjgYMiYTwwus1Y0bkUg2
v9CmaHTokN2yVhhMm5A0gsOEZp51b2kUlJemte9izg7k+d7Nt6xhGSfPAayXfNt2RDgFvRaVTrTV
LGmKuGLTEkzqaPTBy4eCTHq6sHtbTbNItGMM5f3ZQV0XyfPqZqLCCMRxssqlMA9OmnZ5/Q71BGQP
i9U0gOnh48j5OGOqN8TSIQ2Sn71bHTHcOryIXDirWJQInQ1+yJL7G9Swr6v7stuQeqjF0tbve25X
/C16V8DURaMt8UWr1y6vziZSBzy8Vu1G5QYEjuzGh0cV4BRY1IEEiMUZGkjHMzHIi93vVBknCe55
qjNU/3pDVvtrpa9BfKFmD33o5Kiu5/Ihu0lNlo3UoyZxtIZXr9jPeO0gIyT8BkmMIUeaqUnEtzc7
eh0+EzvwQ26BoqFCCx4AbaqPXKkHKQPXnU4pwIq0LWIAW9lJVddH8h2y22Yul02qISyMr1SxP5jQ
Yds/AaF2RNuM73FH/Qn5IMoruDf7y1b5K83pc71lKAyLVOaYR1QcfILOq2hsOIQ86LRacHedSEXb
DxddPgjEXpOpOzQi4MksUFFfB380ARqE8nhioMXftBYMY5I1ouvRTrAJpidJDc29JWZSzqEWXgXc
QCalXfK9hC9OggBnW+6wwUmAeobCcHuCxROLojtvMxBaH8wjdX2D8+vt1qdMsUHi9wyyFkipEAWq
8QxYTIkKz+CkTEcqPZsXPjk+p4ln2piFy+CehNqW2IGnZq43hHVrEYMhKovsxkeaeJeFGnSYutMq
Ri2Ds4II9nJdQZOiuAGCwjq2EvLe71OppGkst/eUBbq1tCOIRs7gy6/7XVFKI31U4EvmHqWfSbPX
WYogDk/pzYYSskgefy+1vDW98TW8fLjzwSwj2A0pJsK3JK/zYT6SMZSMGWAU7jediyiia1KBHuHQ
l2Q3SgvP+KfOq6TnR8eYybujJo5dLwtTdvyWIB8zEOwnr2qU1eZ0NbxvdeNsY0Qjv7/Fpwamh+dM
Q68C4C0xWY3NzRd8AT8CwX1Ykgpwx3yDYAzVotgWlY60uNjoLm3V34Ad5xtEi7+JDdRD99u+rNv3
PHJ55eCAQZzGxGS77yCiFmNVKLofn2InPYdBmJcDNZ4Eymdw+j6WtzUseVQ0lmJEtP9COKDLpVmJ
XNGk1QYq7Gvty+Sk3rY1RykS2665kI0uyeM3EHNKtY3Ub2wZMFj0+pTtaf/zdlRVshMkMKi3IbWK
/uZwQIUoDiQZslKh4LQL76sbNwpnJTmeREheiFHtBS+UAujSQPHfUUP/hS2DjM/U7GrMqJOas6Np
WAUf5mBS7dZXgbUwXrV+jBdq5AupCFuJDH2CefvK2WTUOPHhtA2xpH+Y6EpeZxQ5BcC1+vul8nGZ
dHlit4mFO7rLKLMAcR9SQdrjjj3EPCKrF+P8vrrGyUeXj6d2QWb4muUckzUVWxrxu8YvDcheQ1gN
DuDPPCFyxn7ldVlq7bYoMIGv2AW1LxNbs5Xiighotsh9PRb2K24dvn7GhqgDkzYk1xkNw8xs/ru/
BC4sTAD0TvCDpL2rjN6M1ojPHg7pOK6rPpB5iNA02rSb6SQjYjPknG6Ll8bG+n9iw/gcAzsxiQkb
sdN4T5njHuTg0BWhcym/hk5gXcIqVKHwuFvOgRNul4raivT+uGxTtvYdnr1amIGJ8BY79GrUI206
GmWDb2rONUKaD/nUI2kwXAGgKLWnrGADl/07qyg0V8yE6yYpjwfoLqV72QJm0tXBfjLK2LKvRQUi
cBoQGkkOd6kCX2mPBJQhzyoyolOYxywMiMdvCUfeIv87C/amrlovy3XON+t3jG7bcH4KkPQFUnhk
9YN3Y5v41rQbjeX2fzIzrtCP4oJS/UeWBnKLeF+CS9jNQx7jZLdAjVswm8zZsUZsZ66EaMFlrE3F
iAePZgARqGi9rc+swKzqQpKDwcWhm9lhGGEEPY0x4EWW+7a2wUnRbsoODQjXOqdD1P6xdn5iNfEG
PIOJBS+rjPapuLHAfYSmfFV1fR908e0OaB2mUHMTZh3h2yXS3QcqWzR7D5BfdoR7ERTt7NTIhIgO
EVB2/361a5I0Dywm+jN1X+yGzX813hMwcNGBbtfx8UiFIm0kpnAUOwTuDKcFIvxYMNR72LFMXKG3
lo/ofQFovCwQ+/DxxmhYj4m9F1f908ChkMXyde1PiMAwD/BjxVpkqapeXLds/GDp83PiVmWwzs93
AkWH6JCOdPWdL2M7mZR4a9wrluFdeJh32lmjxZkwQXo5RKPBAgINnW+DrLV51cdwRfq5hnJG556x
GffpD2b1Xmgdls2awqgbpEs2j5sVcBRGknoquPZMQl4PyzH/uPQ81vHVLekJdA7AkHwgKbfnGwKe
l2lsaLfxPf5iklaTFiNFPssjkSkg29fCYFSBJdIq8FRwajYmnVevYVgxLKvRkt1eEfHzvCVKlltj
+aeXp7l/J5LUMTwDTWscHELgQvCBuLUx+qPto5kLDzEoxmNpRdtzguRY2LyKVqJlNq+mSgCwf0iR
XSXew40LDAFNMAicsN3IDyta9kyHVEEVQNphiDk89Vq96i6vrv40PtA70pnQ8oCYm9lKsuSA0fy/
FFpnUlbuInKymRcp5XX82l8/a+NV40HFufxRdcnsfJp2fnPBbdujBaa9e0fSs+lzcOKwn9r4lKHZ
EyuRU+2SU6qvrtjmbwbCGMJ+580eZlBKqpqP8rSLQlJFQMAOJvZDjtnJgHqqohz/CII9vTp8EtT9
SwXNgr0y3ofN5R5eFhKiboU0BN4GkMNXWswJUJvl/KcDOdXp1fABQ31uo6G30qq/uon/AfTzalsC
9SreHRyDa24gB2KRcfnXdkeRsPccNQdsLemUv66Mm4HiC1yJeccN8ekVLUcO74Mbkj08ZMjePUry
MIyaqeOk6KB3CgizLwxkCQ8b3PI0S227KilXSinGiMam1RfMsJXVTJma868+dyKdYFVOtHxA48ln
8WO2dpMitvoW7hJw6x8eaKULASQmD2g7Z7tq3VY+sLPCXvm2OsqHnseR0q7beIwaVLtobpstvHCR
+yyy/mUrVmAxdaib1uDJyKMCWAIywAcJLlVn76U6vt8Yptp5yRmTeaGxCPPe67tAVATX8+E37+t+
Ppxtc/yiPI2xqYiu0euJA/IRilf9QA4bp5wUWHTmutPn0AteegvbXE/OEd0QAoUr5BpzlYZ/P7Pk
AmDBF8CtQpxFOq8TzoHvSgHFDga9Rvu07QM+gacvNER+EVfWsvDEwyL3Slwt8Duy8l6qTS13XJth
o/sI0elv1EjM/X4usUjC4Bd1reapvpJvNKcTU2G+g+7HDWaoDaxwFd6H6+ZHskd/D5xaWFw0e0/B
f+3FLsyonGXltg1/r/gNzy246h4hrNREr5YgnUooZ0mLz6dyzNiLgjuPN35Z8S7A8Dv8hpbo9QTw
N+68GSm7NBmbrvtT5cFN0ImPVotEnySV9/n/jgYiw/KydhQQ8tygW1vlM3fIq45BFOqaQvB4RFuN
6KIrbwTXpUt7tyMywb0nEnJDwxeavkoDtBzJ8K5Ozl2Oin28BXmDUALkQqqqPgTTde44kAvFuh/n
9YhOd5gc5tvDI0PXPxvLHVXTdBpplT5p81HelszVG+ik5XEoAKQ9VKy0YYEJmFmewvmCGOnmfBnq
fgbY2Sc1SNcq6kqC9Y8L5EBNkaILQT+GhRVg62LIJBzdNTKZLi51ucHZxymBaWLm6Va6CygNoGVH
4U0zl+lZIm14gihCbbcq80yBQuK9eKOZNzNkGD7vAlvsoNzV8qjkP4RmBJJfQaX56Ttsh8fJwYxp
ZmfKJnuvHA/30Gwe0cw8DBz81hgu4ZYhkgVcE9N2Y8dJKuMKn3RSCcm6P41T9hpj3+yr0YwUcs4i
Pq2PfNKulsaRKzZaK/8o+/pINitkRPRN5FFMLBli73kDJmk5hVfxW/7pZAl32s4qWTkq56XmmrfC
R3owbUsel/PoNJFSOIto74AlXTUWOHlM6ZOGnS3aG6Pu7LmFoBqVC7KlZPRTnxuQ7iFxUm+UlvG9
oAhZK4e6/gTh3cRkqLuUjJHi9CUNtQoKKjekiFDbz8ttLae0vjpTBrGWaan9lMugEDPx/YjGJf8n
qqHnn3ojjYNHAypxoTjFkhtdoWJ1oqmk/DSDU1tMZIp4zQrChVDfTh7yDN17hkPo4QepaJPG5TzA
3KuxmxXVSs3lcnyixdGX1mvZ7XXD1I0xzqWNH8ItFKXPAieRzR9cpgsnRNkKOA20DOEL5RQEy5FG
IFwqkQPx5nOPzlzrDXJlNRkb3EJvstyzuhLtmj3z1aBWUh4Xk1BA3OTPET2KhuTO25IYJbTmGIyi
NC/BqtNCI6pQSoLYoTq+yer8Kc2xyy52BpKWSCWD1Se1fgd7CxG55SIAKMYQj5B5M3Otw/HWnnu4
TVXcJHE77BOZVT32+ZHfPjLIsAnmzj0IcQA7d7ybnDd632NY443JZcPWEQrhAMoMzLfh4EkZXU59
RJNIhuVAnamc3TyDokoy3rkoIYzjBrSUUL/9WmlS19SQdxrm3cRKtMw3CWjWF6qmcOR5PZ+PjsHf
o2tfHVDGL6pTdtSwgppQVWUmO+neJdX96UYrtJYEBO++/K1po6+1k25BEwfz0sOVZ/SWFheMq2sJ
hJLEorXktoJCplPolEdBvfw27ZLv9AsoHVJfKIhqK82dFuP8Zme07SGrKZ2aIcQw9eAIV8Hw2DYS
6smBlSuLWSb/mCs4+gFRpYJ6Zl1W+aU+Bfu6Rb5KwLCDlB6NYRmoyqqkRnlO8wS3S35wBtT9/5nU
C8X93zGebXfIJvP9O4wY1pEzKpeCcft2lQ5azwszZYqwaXaD3AW1Ih3l8dwG2LLdGMAR7mX6DJW7
ZlTKqEvTnzp/G2OHjacNtH1lmHxKQ6LOEV+3zxsiRUx/FyBFzv0i02t36+oALzC0/tYPh/FFqV4f
6jx7F/M7GTwGmrjntIT0790WgykWT28gwI9PMa7X90fjhrfwXWAihCD9kCOOgt96DpDvGn4S8x5W
X4QubN43uNjoW9gbzfDbnfJHl5yqluwgQxm1c9dnbjWd3My5G2JWsOB4EcBgjunXZM3dcPhhPdrl
J1J1oqWb2ZkpnutwCH5wyQWlDG2swqjCnhxy3CrH7dpE9iOvqlV9orE8LhAepMCpFi9SqC3zS1lR
FtNb8LtopcXTJzOyzGvz0Ke3ZMLzVwG+j1Y1bP0iGCr20rSjmchIu9tBRk9moKP20Ea5XGA1BVNX
2e+ZhM+m+O40/lBkrAZCdBckNM8Vrb1JMoT7jKu0U61degSdu4EcgXEourpclAuetb8opBXlsewM
PZtNqp9kpfmRj7Gw1yNmH2kysCACfS6gjQ/KLfqFfEIKBFB+yTPrEjrK+2hUhZgG1XhuAWDqWtQa
0DYOtejjoNruU8/PyL7mdhZXV95zrAd60nhmM9bRhG1G8D3bFXEmd/JzUxLJRFYCLmECB5I/KRMC
0jdzgzqPF2DrIfD33+XosV7rueTfj5GeeUP/GlXkOAd2vHH41SDVuPeljd3AgrJk6EJPfxIqRAIY
v0vNU/75mbU0eA+W9bDnk9SsxJyLZ0UfK4S+Co2+tjg738pPDHoi8LR4l3G+EMNMR0RPZah0Hw9v
JWzgiBGH/DqsUed8L/gusqn8VCs+D1sYnpMDnnvF96KqmOAAgo5769aX8N/gH2DdX77/BxBXZws3
dnQKuXAaT3Ew1JiHqmUdztXKOBcj5Q4i3GZIWN4vqsT/KTtDxWO93NiX9+zyZs7xEcuER0j9kg17
aFXDkNv7yEkxw4UMhxL+cSl52GVrKaXtLVVK4DXMSNRSNnP2TaOplkYgyjPtggrd6+6fNK27Z1Bh
eivLqKiAIUKMKfR3Qhd/d5tWe4mmsfZiT3vqTegf3j/I2CCjUpFN4tEsaTLwHRbY15SqRnaaaxR/
axqTPfRWoVGnen92edoFvzrym/z/sTQK4f9vIHYgupbMsCH7cWiSyXtwyu6VcHeLrhBOfZbgZXND
90KwMilClSWpsLHHod37zGgtq1+w+ABRRgJik68plRAYJ+JvVCwwOIRKKm1/bzPoxPL3PQzhN9SK
F+DnMgOXIn38NyL1xUwjiF0dhHpbm3VhGkNO9Lb90s1QUCruDYjbDkChC8IU5ZLlL7AUJ1DtKie+
wq/Rmwa5sJRndTONPQJIv2QC+6Fow4gXcJ8dbVOedf09JU1TFO7HwSQaKobcwM/sDbbpNmf5al/x
ijsQvn1aeqWSsIzxdyyeIfeULRpPLhXqTMRyilr6JDXmk714Q+fQw0XdtK63mwkRhv3zVID5F3sh
OenenitgU5jmO6LHoR0lIXo8i62ZbZwNHz2UnDB8QOlysNGcoYA5jOSth5kYwjfiXpewkpmVXgwA
zGPQQV14U1xJ2cxTGF82Z0Or6jbuhDm9hmYpKykLYGPvh1gL2BiKMmJHtrvs4rMfelcU4QOg0Cqo
s85WCXww9351oRxjBWNtVH6hCwZTO8iziroH1W50OJvW+vZ5XAiyBkRrHZmKamv9fJ/FuyZUo8z+
mxUFsEgdp2h+5xVugapbW2wZixX6roO/MIWC0Z4rPvynaGYX26+4nFjUQw4XnqRrv/QBk8viBZJW
ULL8rSO4TmZgUdkofPtqlPj1nviB8NfGIlfDBkq5UBBGrX4ypbtm9JmUFi9ltmWrw5g1r0jcpAoz
Dtp2Sdoi8Hd1hfjxPPreGDAmyXheXbRhMLlmCmo/FVKpTaoiuKBGy4lw/8S7xRciAfv8jtBgA2wm
XowLrxZeKy77OfPyYv1sG4F8hI+aQqWss+IRxxu8tRZQwFy8/YWXMBFJ12TYLyUqep7V0poLrZ5R
QMpMLhYEGNhPfc+KijiB6NfVbNCfx7T5H1ur6zd9rvtaXChuyJ9P8Nb1DWPkjA00Qm2lCHMIwIcz
Ytk9TIt34gUC9pqUfBUN+ogaLafxk6A2BPirOhDuBu+B5/ONEj5gl+okEkfb68hNfXStv+aXiG6O
4oXVt6p1L+giNzM0VfIysAvFFxbL//99ciiPhyIFwH1TFyhP2vsmZsAZCzN09ydcA/m6helS+gIR
JuVsR+GpnVyqzdGjvM8+1hgYPR2urZM4YS725VwuFQx3uqaAZt6xxP48F0+I6PHiPvK52NKgpuO+
r5B55+V0PBHCzLghjP0hHCmCSInviyKtTeFCepcrxntc6S7MZTxpg9qi0zQb+PFcjMHIw3AOo3pw
HI1a9Z5GA5AUhGIWpiEgGOx0wb+Agwm9kH//I+bBJZ8Na538I4O9wtLNRMscnFDShs7pB5ivDeFZ
Q00lhjZeXzoSuyF/sEGTIcluW8RxdU8oJwxxrkuLb5qV+XhG8oJ81jetF0hJ7pmL4yFg0MJ3pED7
qC2talAraszjXH58N8drHj4gSFW73L0lreaTatfoqD9yyrmzLJJzkZWXKL6wfzJwKUBxp7Z7y+bB
iklz0sn5t/lR76H3lh0x7AEvOohd6w3J+JTmuH+4jfGJNncIq3H6QEMTk5/xy6h3F7e8XB9EPJYX
20OR0osH4daQbmSPNtPpZ8SB12Ep2KoHC3RuaEUtVWgrinVD4tJhqKrg5HY47nwP+/rArOr5vVbW
LN1/PUDzNVJHTDtoAYUsgBTMSZ1YumX/UkFqJ2FTvx81XbMmTV7PTLNLP6wAOHYN+HzHDwJ/UP+G
Lw4+vji7P5ByOP623sAXCo/FlDSC9g6oA2wuE3Q4kNDsDLPE2cz69OGUZqKa7j928qJxnWe6CCwi
zmLZ/6Xh430zuikvyWgn9FEG+WVkT1WTCjHe+9k0N43+mBL3w3D7lCzujwqXDK1jbalffOUE6UQc
6U6TiYcZ6kJSU751ed9korHrg70TA1Nr/3YKm6C1JSJai+W58rMQO+qTmt2BJ69nfIll/GCziD/3
lWDJhtal4xr0HejPmVwYX7hBotr3SXvhmGZHOOGRY01lJfZ6G9hI9l2GDwu+QeUzqfwKC4DOpsBC
lEEVNCGdcOLChisFn31rblQpXzeUwM5/qaTSmPX21+0xJRZztMVRij2+6OpBKcAcfbxCVcxCtZ4A
QfLsr0OUAkx1A/sna1UKfBnc7OLETNIzxrBzUTOFQ2FnJNI8fqP7AmaZbFN0PXtDzaFDKZ7i+0us
QZSclUFgNcWbHLJ9pKhXqiiBhnSIHoqYI/K/CJkcMTTnTXQzsfXLKfDyRfKU/VpLafnn8y4Q8X6/
ebrG393zHJVa60LyBb2P21Y1YVHnPPp6j+lnP99/msPF0CJ4BlLTLuczNtdKCLxLa/ZdDJgVXizU
YCjvL9CJfGCSR4XJkiwidbeEtys8VYNAfVbofTi/vxDbTJZrJIM7xFQUny2OoolQ3AoEEG6mkh14
9HB1EFZDRYR2qVkuxhAn3DGkNL5sz8sQCfCMUQ+bBHvXiYHs7bVy/AdzOZ+YVprezXAzojzP3mOY
eTSOY+uNtxKBWtXuTujt/W51prM9iw7PvmYEgwQV2FLZBEdM5Voht98kt6pm7zi55Anq/XvAzXAJ
dR/uTlHk+fZqSU0exN6qEuXlG3LFcgrcEPaxJYhQ4IvlL39QEkQX/0LYtG2FAoNEABWjVR04yBqc
JWyqO2LAsSgOx/mAhNEeA2KAYSQCh/fo069+2VmsUHD+vmKHZfZpHvKTirlMUjMG+u17evA6EJSs
HZPAD2/vme7F3vu+oWcdR/Q4BrTlw6G4INebcypFbT3twQ29TYItDd5iLf2VmZs+k6amw8s6HEEQ
JW9rrp3YpInAagL7IMiETsRSYygvjH/g+AuMUcQHhcv46OobjBkGy5kdkP4FhRNyaWsQ8H12DP04
vuesKGnb+fG89Mhlt2HYGSgV+mLgpZIyiiGtpmRi/f9k4P80kV9whrILfX6BaCerT6RE0IiGjROL
m7S/pArzMNzjG+NaWmaB8Ic8EP4hjjmvvKVVIVk/KOMCj5WBA5nCwSam5in+UI3jWU919Et10TZ0
EgDhLqBJDiWsJJW8CDbgFAFaLHPrNQWvZTg2UCrgRRVLSB2Zr6pwxlYEvCP6XUcvQtCoPjc010RK
YECMydQ0LqLfVUzuMbyXBy9GNubppfS4U32eHZjVm0R02yGfuDLOBn7K+5kQTt4Tgrkwi9J3ox1C
Pqo3htUf5NCEorRIe32VsCpdszXYSa+su7QV8E2ZNfwtaGWfZlX9+bX41OG7uyYf/Tc/Ulq97xFO
MSWtr2u7MpaDZRhJZRC7D8Tk8MhoK56fY5gWM9F9Gtz2f6YvzssU7XTvCYZSUaGuZp5wt49C9OJS
WvxH3C7mPDncGn9Guu/U+f9nOXltsUVpx45SsumAwstwutW8eDv9LSJGHweZIjD40HV5UUHDmgFj
S4FatcXFSaF9+G05apja1/bnm9OmW/3gh+tT1FeZxGXSsDs4KOH2oKLovLrpPi6yNwuZigjf2yuA
VRFTf+vYf0ijWT6+Uk/G1qEsmJMc7AUxAC5lKHqUYagS/5qep+nfqlQBmrGX3eOMJ19QVu0TdX6G
8BetzPuDMHtDzWB8nHEeOvQnirVM3fwuNGv8ysKkMzP6ZXG87LQ2h0RMctaggrN1I9+nSZsHLlGC
TXS0MJsfwlWP2+JzdGkTi+fZuAtRifCd3oBaezHwwCJFj3HrFt76r2ynSMYDGIH0VQCY5goaMbIo
lyS1EzyztKVIfhRUqW64ru2cmb/Jw/jTOlnKsbhzm/MXyPpgV/bU/GbcY1fpQhw7bB96o7f/tHhL
bXb90o1EKOCdR2JYxTVSbmx3zbwjmbPinL5hTH+NxGn8cPscNNyw+zZI2PVybFpYm8PfZOgLbfTt
Ui5ZbIrhgfRE5Fw9CzuuCqa4fxdJNkMK+pkHoGNxWXILG4FWx1spNxuQ1TybUTlkqccQLhMzmfRR
do+Ua1heLsNTtx5qYZgKIUqJDrbjfZ5TRibBy4csSt9NrX39wGYzO9BtiwNesQOc5wHk+0y3rt6d
3uktC+/ATwOEJKma1PxARzEzk2HeHO83WX8upgSbVPtKwLt+V8S3h24RN2UB09kg/MDFMLOxJzfE
4FvgqbnYODz3alNYDAnzmIBiIjI4DmzKF4FjUohyOxOUYby7mICjFXAVPDgCeiLamA2m/Jmv12vY
1GNcvtE4kWe+TgrmifpLY41ER5v6LrEFLLOPw0Tg+stIl6fvwycBEKeMN7cfLhWtqS2KMwtlZXyC
dvPT/nSayXXgtIqi8ocwl25wbFyzMrzO3NKStqMizw5vatVB6q6acUe7nNlSE6NWfukXDngHF/j3
m+DeG6q1sc+vXyQrKasDRMCYfkbG34rtU8eyqbTLgKy/mniBU6pMsgdV9OMjKhlCupIwKu0jfQN1
/tpmqYjx/o3kn2LP4qjnyO/nIUQD+7UnByaYdGP8zSn2AYOGZqUukfmywzX3cmyGmGy9h0jf2mkV
K6N0ywPfqO8CMna2IT0BEaHki+R7RAleCwlrDFi0NlKcgiZLvoTIYiIMQV3YunOGNLLGRWfGmJTA
magT0Bf4RDaGbt36pfAtwv4k6ITTpeBSCB0tlE5p4CF708HAYL68Fn3Lh8Kv5hfEsPMmVwgB+4u1
BEmf+JaAjAx/hUEU2lPW5gxhgOHMdCzGJYhEuQOCYpBbCA05aWaIF7to55UjEv8gTd9eGmURi5ox
cht/5xyW7UTqg9bUfBh7F+ZDvmV9KTSycA2x8shooVQA12Nxn/a8FBIdMsilTuvxORPtscqTJcDB
wZxuT9e1aVsnCfrM9VAnBqAwIBSW9VctIwxl4DCAKNCCYkfIoXG2+yUxWVo9wvRwEjmc+KVn2Sf0
M3Cz5brtD7OusW3lOhdwnU14bC5b7CeFouA1of64Xz89TLkK1BrtB30SCwiBY6m7fWD6iMbju3/z
LkxanFdiJAO1acC/5KWCWanGVqC1eGkA3W7ndVS0mluenIL8aprhP1WxvFJpAQgfKYXmbzs8ISI6
BqTZVoxn4T7pnSUPYKf20ldhPhNdr8CrW/xCyCdeR7q5rVGI3fENC64fylGcGdo1wRqimYCY7BdV
fshCHVI2EXG/hnPEqenEfqqhWjd4pGZEploQ2HMToFE7DoGqJExBpbnl1J/q8CnpD0r5Ys50L0yo
TbOOb9TmfVSxtsq3nP0HADAaaRguwSF6dSHNRZKdo6TZtG0DUYEM4J8BLMuq9W928hFqBFIO42C8
Bo29n9wTr9dq1MwfjMl7rF26En87ScFWpE4bt3GUXdwtk8drSR31NkKSJnnBtXTfzUTI33QRlw0g
UOvi6bBH3ytyXZa7+O95HrAJNLiG0tTY5xLjgSoRY8A0F2Zf2BE0crrWdKupDLZJ1FS98g8PbCtI
yhkwtT4UZYil81vDT80GTZACdGuyxzoJA80Iu5WTWd6+1qkFEt1qQvpxEesnfwxr/JK4NooUw5wQ
naWp1POIbUEp0WzQbaiCZ5VKizchXZM4GOisQzxvQEYWVGbInw0Z1kl6JMBJqCPZlAJBfK8WhZLw
pXGINsG/VSuKpCqB3lmZ1FYyR/xGL9DNMS6zrUcHX2BO0Ad7cKa4GSp8pRfsDkaOmtfR8T+0SkPR
//0ba1Fhv5EqXFERg8ffsLs+UiuQxn4ovkJOgxU6/OptS27M1EDPL9BNm9SjXGnq7d3FZcCoARqJ
OWEDNWhC9QQ02YUDPGCRLhspU+vPZ5iu8yQVV9zKeH+PAJNau/6wutWA+JohAbjXgl/ir8y55cf8
QvLZXcNKkDouSyXOiYLYyxfRuElyBzfR7J4IWkB9iPbwPhWTPXIqvNInFUj2ph5eW8HVPbBtrb+S
Q3+attk10V4hFVVfK+G+6yUd2TsgkiFnwPd9MIx/tOidxKeP/Jpol8qgxW0itnv/T88w1KCrV1Kz
jH4QiLbgHJC7emc4Ycr96rs5lB3BsiO9n4YYuuK6zzo8ai23YynATIwVuleQLGlo5vDwSkps8aom
otkG23MdwQk2vF5zKzZ6tKITTQuFLKrL5cLX8SuQI2rCB3KzfDpB/IQmXbOHWNxISdtYpB71aXyw
ovR+MpVmwG6nAoRrWo40KyDvNtmm2xobFLpLqEbJkSgwVAmc2n/GidNW+nFlQfRgv5/rTUQ3UI5e
k/z4ep7x8XuuQagUTbfTR16VZUF8hX3ye4/MgzsjuA9dlE3y3F0CbQHnJHFbCKWAn+vCL/sKMBx3
HvjOfTUnTe9jPGZfOkq/R9rJSf3zQWiiCHH7ScyoihHdHpbWU8VcZ71AEJXsky/CoEV/a7m13Stt
/Zm+nk6i5O+D6hzHGJJKJ3nEUPpFwCQIm+OPm9Lzt6g2W4deofMpPflkWj/nM9GXBD9yXIIjWcAF
Rpk/gSxNZtTwxRv4Qd9Oth/YMRKGhV+1O8vsufdt42KcKfBi3k0G5+9oFST47vfl5ufGUPeMAXo4
55wclfyl9GiHPsedgTxPFjSycqPcIJTLw7Hl6OP8U+vPRe/6fQTJ/f+s7nhWmay0yMP69tfaRgOG
QU6XuSSG308x4eTXJ/kYrbUP6fUAf5I9FkbK+DaRYmC4+nAb+3+EkIql//gNsxfLQH+HiY2PJGTC
WPGclvrvept6AHuhH8k9k7gZKWQO0px6zeuq2Pr2031EET5DiWi+v6Jzt0SQAV5qqM5V+DSQmPGl
V3QlkWpz0GH/N9QMsEt57TEL3E4h4SVX+4QaqdLlF/KB6tXaw5A5sPYathuf6fDh/+2JAo6GllWI
FIwaarLJpL7npZ4B3IfP2jOuDAgwxZEzu566uTIa0yCp8B2swUufNtbO5KWZt8T8avSMFDObbCSm
ntFcOdxtSNyX1H9Mv5A2WlLTdrNdvtpqDAYwhbSKjLrf8yFHam3YsNM4LjHfZckO2jKlbHi8igQf
ZhdbUxEo7Irp0B3O/Sj0f+6E6nzx/cHQEZCg9aeCL4Hlf8e+jqrA/4qOG3PJfQc5gp/vKKOS8DSs
5OuekboK7cg2ThHWiPL7UANkGifuRsx9zcRIScanE05oEv1myaqrGKiSGUa3ezZn/I9AyrMm8CFN
10hGMTUHptsgirJUG6uKr1WV0x5c8IjwH4+eBgx1yH5xIXZDNXiQQDHA9LecsN0uwY3wK/McgcOX
eeguZao5k8yGhr2M/pFQSvgRurl+vxElWanlcYcz0FpWoyRhZGM0JV7kHvsgwXcQttOpOz3MOTrn
z8cDR9fgS5/1NLcF/d78KUrWHIaG6GEiywcKpO74oke+mIvLYPTDumkFIBoLq/03tigEY3QV6zcX
s1Yrqnw/goJb6+6frZOm8Ag90jT7HPIMHCbP/P3xffZjAgMRIdRNY098XfiTcdLg3F+kIjQKIDsD
cUjiaWCvY+Y5HV9rL/GaZNMsc5e3loPeuJ//Yo3RPxUq+Fx1t6SmxqH3OwGlSUNpLK5x030EMkOs
WQkFbJwzh9pv5Gal7OuDr+5ttaUE1OoV+/s5moXvgwgHjXzctFxkX0LY97aP+hKbDNw7WQ++1k/h
kLVuf0ArSZzM6rT8tCsMzvBWccHcHUOqCgQnTprvNb6Wft2PNJgbscDj74R904t45Pog/av8Yrb2
uQl1x8yStOZfWfgpv++KhYRCyRweXXI2buG/4vz1WZ/GB/hC1LZj93254lxgg4uVF9Esk/XKM+6e
MBze3XW3cwxhPOOTH5RpBnfWJDx246aRIBqtAzHTw3v999mW/0ZdoS46iM6KcW/Z8TKQsUQbHapV
5sakYtjTDN6Gm0dRLIiaD+oWG4vbL46FEGwLC9eOKz4r8RuugfM3kx4z+jRY5NpbMZjG6GGyYrCF
mlJNlZ0tjrx8ivtQXa2hqU9jhm8aIQWZaYAEVdLufBQ+mgQAmtJFJTQDZchOA4UT53tbaZM01Hk5
cneI5UbSZby2Y+zqyHFIghXHh1WRjdORybKhahW8qbQVjZB185zaYZVxZdYPg6XeSrgmsleDg+Vg
E3zTfW9Oj/4r0lAN+MkpZEyazmyE5O44iXuXqrGRv0kQhXLUoy2UfRoHBqRo3eESvGnBOCN4BP+/
7cRrQdxg5JGykrh4e6PYB5TifKyfmD6f3RyE6hphu9sZC72V6V2L+0uU60reCsHs07/a/tMyzHWk
8M8zKQbh4x4J3LnL0dLK0Bvc35lbftq+OhiagJDCEt7bAze4Tk2QpqzoJJDBeoPBHGAb+5Y4/RLx
HkTjgjJjILr/JKcFuP6fvrS3JQQzODqEF5OHDrs6hTpu2tlVvEodiB2UxRjEy3AO+GjTLIMhtRI+
dJ6pPnkTpHe/xwFIRUwa96EzE0gAc1C32mhphGtnjqnLtKALDW4o3+6G7iHbgwlP6I8dNn9BtqMf
wuXpOLxZ/qYnyFP4Q27SCQ1JnbKR+NpfRLHUCulT7cHCAXQo8FRtTRKd4m2IiDFm+7rF5yxJ+iPa
2m+NOq4KdGDHird9osrfXD1YlpQkBWOiXl1X6IbwRYQroXQt5TYJSAdrxl3qfEl4RvfCGrJuxi1b
0wWkT5UIJo5L0fG3ZiIP7WK1FHXx+90LrxWYOWyD83//2fAXO4f5Tm2qfu0S/VOPqJpFd12KU5CB
nmKWL6Nge4PVHiy9u0yvV0a0awvcZju20jW3UzJhgwmLrv2EnfO4m3jHMg+59z6DZbWL58Z/rxPx
7luZjMmkCJ+LYH5lssR6GXe+BPToF6RXAKJoihODEzElxHwwB2UCym/li/X5SBFE/H4FFyQKYGvC
2cQ2WLFuwHE+nWMw4ZQX7Bvz9xwaERQiDzyummNiiiljYHYHazI6kznBoQYqtpjwyt/zPz1BoXwz
rWe+pxX+0yTwPzzq9C8+XDAjFv9Pcu5CGWjNuBV6zbAq+g+sCeGC5JyN17hc9Y0ZsV07XoubYzG4
zlM3MqS8rTOqnMuAO+zGWga0nhjrlzwheNFIwKR4dAha3Ow9VuB1vZORU6Lf4h/cMUwGP0jv87gB
FLS+XhmdwG4ME3aOLJBO/vNxya9KhamnQ6RkY6kfqGIkebWRcOCouyF4KTXg6FPvCSXRNyOkFP1G
QXJmAm/sGuQOIQQR7XXGaTO3zEwlNLAUIo0K+uqeqrEcT8XUFQQIChepc7GMLtgXylVC6YcQaBkK
885tY2E++dj6DuEfwJgdTxs2Ejf8tNszXByTFaiyQdcebnykdb2nnWtwuoMy+mNmNy7t5cN5Nzpk
jhzvlqrB9xMP8cmDqQSYaTXpzXXmLbC0udGAYC8hy7VQJZm3GOW6zMX0H/5G7BptX7mCMbhATNJo
ew+2dbj0ThpwVzN6djzg4Z5s1euLuogSiO9VzC43ASjWIUxwrYtrzFrvj2uja6sla3FiGv3vvaAX
3aLJy4tEaFA5Bv9lMxZ8faIgQdcmAmC5f+l4iP09VUiMqj/wm4wdQRJ5WX1mm0NTERSHrgByB58L
gl639ZtTfcQCBokKfg0ICln9PXIFYVhRlNdjhRc96lFSExpmmKc4wrwvF2Yyl9fkPvVbr1R+wQS2
I2p6niVJrTzelLkjIOfasdTYumAEarVOTBeG+PxJmW9nrR4HxVq7pxDYWjPA7kXhRrKUdWJrQJI1
p6HfM9v/1nS8968RkTz5XPSQ7sZqlXJA8cMV0TrpzLcnfRn9YaCZyDh+MqUkX8HI6LFznL6F/Au5
Mddo102NiVWGwN+bn47ayjXN6YGZgeb42dzQv0BNttb2lVNYe6+B3XpxQHqKU+Qd1kYmOSaSmQT4
lP6Zp/dWYTG756OZqL0cKw1s01PwwcdBVVQ44CUUBpV5uOFEgdobS2q04c3CVZT/annkMeGY1dML
8/7KNp5gIn6JrVuNTehuxu4rsMVTk1DyOcgbJzp5xrMULq2Z5mnskspPNtac05Ffdjm1RP22SKfe
aoVRrxo96tI4S60LvGim+YhUxYyb7/ogcPWRjTu2K9oR7ubIHakQ0Ru38HUA/dIW1FiucG+VMBwz
they8gIdAGKo0TtmExYTr+pI3eq+M5dmha+k3hh6nMTNiU0UxSMvraTeZ/47dZjiXsbzIPzk+UkD
ei3WMGLqYyf8CilW+AUNlZWkbyNiDOF3E8BbjHXANZpAva42dZKp87rofvUe+8G0/ssQ4C0SDVap
hJQEO1w0kU6KXby12dnB55M+siBBQEVQEWyL9MSQ8JsImUaHNKAVivvD8mfKVu9owkC7DYin53H3
UP9wbnbPXXocPjIuCtTaNPeHr6aXjDbyf7lINRlMovbOo3Zc0wgmqNDLKc28adXOeN5YFyyk384j
IOV5kbEFfeM78GCPioPWUatHSMN1YgPKsHwKA1cZzVas6x06hHwMGpwuiO4X4OQ+STfDlh/qrx3o
jLC8q/03dVIHW4rKRLE6ctIetZmLxJisyAjw6cse9y/47wJR5SKAnDaEKst0gzTPMIT+PmSvYhlI
rnUFKm57nL9W182aoUvNguZeY0/AFhSP19Uio88DKnQ/bKGYYnwR0zwetdiMWgpYWXMz0nxHBImB
V6v5d8zn96JBmVgBQniAVoJEQHDI426tBgSlr/CsUYphL0ywM7YLcGiS9X2u/jpY5A+2YAcO3qRz
AE2EmumRtt9sKTX8LTu645jJ8FW3iVGK+9rP4YnsUaAqqzrkiGe3Ojjmhr/irlqS+q29wHARhC7+
k04Hm+5kw/pXW6xZTBtpL6lPb0dp6cCe87AGpBhrfKgkQQe/xR9XG53JB84IxUo0he3oO9s/CHm3
fAnUnUqKcwVWAFNoNcBmO0VIRnCV8FPFs9SCilbAZZZ/KzxCho7YPtMpKtnFXfi6DF30TbZE5Rj/
tpgE1cW8ptZ2hJ2lcTQU+TYSKpbLDULr/Lq9LlDkgIKShFLG4aAmVczNyhoM8cEh27Lf9RXQX9yd
ggzs0/MDfhgWvFqMhwHadbKZlIYLq/zOhTpSRmg9eOKTPU0OCI1DdOKa/zJM530uSCAZ6nZT6jKf
6CwPA+vVCes1Q3DVBs3iJQ4iBQfPXUh8a2y5H7NrG+E79RgkyZW2PjoYjSbYiKbriPoRJdEBxL96
vv72gBQbXvep6VnOdIed6+fahg70h8VHTwBieGI5zuzKVh+EnNopbj6o7JHZlI2sZ2BCMQ1rBEho
lDKmqBYc9gmX8Mexz1NZixIDDzIzqwMyIZ51UmFvnJbWTKoh0Bz5BXJjzsRS6Gz4wFLSuZR3wCzu
MGIOGFdv5oZBsf6AJTNUJ4SIhkD6mTpC9CaMMj7UxHAeZJEa/pjP8esGdFdjrna4zSz4v0DxrYbH
XJwUdPCBVIrBVFR3fKdYTVCy2Jo9fSkHn7K9k3xbdsou/4ekhfAd9t+z4gShDBevibGzFHYa3pvY
xJPOmd33sFleAFm7X1E9W92YLLtzuepZHtvauK6oFbMXxFYVCJs7JVGBJ00laJpCPJgUVesqYIMz
piKDXvb9GgR5JY3wfYWAzW0O02PwNieWtinfsxL2fZLiwdM76P+fBNoeWy2x6SBFp3MaKJY0cvBL
f8SjZluGeGRTQtLTeV6rYEh78FVGE0k4gl7249xR+eqqj4LeDDjHSUTwve/hWVeHCm76fvQZqke4
NcS8KcqvFetjN6QeMEXoOfcZs/wc/bGXe5yR90uJIeBAs5Y+xaE4764mG62lST0VUUQnkoVvlY5s
isYCIo2TAVVDAYOsrB6Jzsn1+0c0DoEjsOEsEIq8gi9RsEysQ9kL9l7bWMXkLXkSXjD3DC5WPNla
YZsGE/0kvHlsDM4QepqAJ6zW39x5G/UCkeh/GMStdBrwFSU54qiyaiBac698JCcsLo06J0HUHeSh
j5MC6GVnqV0wu8P3HjY30ttZnED3VeAqG8qIgSxobaUxjVHLxtD40LnrzFKJ+MuNMbV5MF6RPkGi
DYKhVrhu/9BRzLwFlmyIbB37JXfjKcEbAjuZ3hhkIFC5+mqVyB9mGnAP99jgfgR8lObdVlQF6Z7v
JW49ZKGHyxFAVv7wuSydRcPI7uW+XNwUOVXzULlTygF+acbtUV4718QSUJEavhTeuU/FeaqhHOOC
4b9SdV7jYNQ6uIT05+DiLeEVXwR4TBt7oUnxTWTkYvqh4BwjtwwQmvpxYOTXGU+2MiH7EWu4tegk
F5aMsjahH3lbWvhKGo6KnQ+YGFcllnLiwgYR1XwrEeMMQqEJxImEU0XLLI5cri0br4CiGUccF1ft
h1eirqdbcC0pNB/Q00PgREy9t9MW0DCp+M4tiduGxg0kZecjf4jKCpk/YcwUepA72XqvyRuWhaP6
abKGNKomroKfdDoFCjfRpAStmNR99y/6k61n9B3QFDNSKZ3lyEnp4U+NN5bZht75H9+YYuiHk3X+
fYKTjq3kN78gPQH7Q77CzNtiRSa4TCc2p9xXqE94tp0+Era1Qahf+xHGmp717zQqIA9sRiwkIlAh
M2DlYXIh1P2xBsLQ54TRwVJtPtd2Ic2K2JfnxtCsu4qQ6hfZFA+AMTh1viUF1dhq6WdZaPqXBA9n
7cLocJcZ2b7L1r9w+/e5XXIDGLswEdz1w7d/+C2W44YnH741ogZYiE2kmy7+0qpWt+au7IEWZvlY
GZlQvp+RI+IJtH9SWzHxfdjqjl16Sz8GsFwplb56wy0k5k5nqCIgGwuwWrJtIXNbZ9+Knw9Wf+cI
K3ySFxmwVB5gBi7VuazMR9dlhBp/ehj2WQwE6w8gUF0z7l7JoFrvEjzUFFTkDAqOSomTKAd/9xl3
lafridxgxVao389MwjsMXRur/0WNuNTUJT+ECx79T9HECQkLCKSN4UK9RVywuW48e9akXkMF1ipP
VR5PH595KEGkeqS0lNdK179DZmUhFRCqZFUX0Jlw32hIbSpv91fyLEC8MqYuq1um2E8va/THJ+jl
aa/eu8t00vuVq5rcda6b9/CxzSbznXIN3WfbcD7WyJsdemaj4XNqmUrhF/beOGzRpV7IK8gtcVUO
BlNQ0tszTjOIC0wXsxEww9/9EERwliBEUGD9dTSmfqoA3KypxMFR4JMzQm/xCORSc45X7KAv2G91
iydxDU8l7Dcad3yG51Hw++850oIRIIecaXFVDh0qW/HyUcw8d+kEvQO+pzfhGxSNCtkClV2PoLH6
KIoANI2ELOGsokMBK83TqKmX2TTzYtAY6lQAqChllObYiMBVH0V+MDUE9xrrjVSbFXJykpWK0tny
vdlpnVi3IU71/wIOMbuDPZtFZrKT8MbuGyxS1+ywWJT+X0QOWHjIq5oJgWvnrxmJQKvotKpdHn4v
dbyyLMobsVucnD3feUDlOuvAmlvzhRWmPel6V5MbfOV9VBMlB+GRxUqrO232m0MuScXiUoHOoOQn
K8a7VtdD9RGO38jQiKWlwmaJ2c94LB5EhOUwFSttgOffAUWVpyP4I4xpU9CJJUyc6i4/hAriiMJE
8eZEfLIjg25GNOy0fe7bgUpMyWPch4//7o+X0HvpxkuWSbAwPbEG28Tv2wVIa9H4kGKAsVFHpv3w
urRM9SCPcaw1Wn6OzmGWGjFHh79wYuJVSepCwfwLbXBkbg4xyoz1nphZNCXwwzaWITPLxN/BTF9f
tj5DGShvFp1Cae4R9afK9jMc+Z2fc7XkiAoj+2BO3qeJPRf1/M+U2d/EnFBahJkamonf6TXLllfe
MEqM8zgjc7b6mJwaPQdfxN1Pn27CdfOPXKlGGudFvyT8sg3h8r9a8J7DnOnNhcDUqNTYi9ayY9Ex
A7dRSCc+XbT5eawaOjipqk556c3H/kR9zDk9Co5vrCn18sy78vOig9h+gybjhKJubh/ZUEHJ4ESx
HWvdtUDphMRU+3bAS/7BtXHJ59oURGkSJwDuTPCbH/STXTrgMNAwt60KMSdEyjV618a+IDqe8pmt
pzAwDVx7L70cbkhmpaXywcBz7mOXJSxedW+sJVnI2b5WsW9f/5HxUGRw4llXbdNGlNdYws4cIp/Q
mfF8wWUSs+LgrxKZPvS4ETw7+v0WXtNgxeO2J3M3+0RdJOw7BKNq5QAAF4vjlXp5FUydRplhlywP
9JfKr5yNZABFAnfjb1JSgs/W8ATVoiZePFo0sTPFRDo4fW7VX8PNRjgOpSX1rAyKkKc0um7/af2X
K8pml+assv2bB+s90I4BVvNAx/SbNDXL60pgev3ZFQC/uAHxyhq2lV8lw0bdEI/36c67ZCKH1Cek
IRALcunDUKXVWMkf2W3KhL+49Gcj0BS++y0/WiR9te/Sx2lJt3axnvko3PDUzuOe80yX1zHaDs8t
XoJBSYoa+UWOM1Qj7iHed1qFG00SZZ1rv+S9wUaXOINjYSJgAWd8+rqXvl008KfUrveyi+8C5blM
GyEGPqMOXPJQwG6GVcSMdKlBExMFkvBqsi9srkY/gPXcSGvDf73zpdxPE2/x0Qh7OkzpzlqjeFDp
MxRIYHq57DGWlvwb2jkW6g/O2Or/dgpkCmSIE7/6jQLEyeG+FaATO/QuxTVHLAPTJlgTfWYfW+87
Flk7/17+9R40R+yhMBVfY94LSlEzOJjn7MZ6UM6NfX74RWrEXZUZUkJDV1jPeLwSRoYcfO71oTbn
VGT8apxrmG4QPBB9Cp144mq4yDLgh51HuWMjgGYi7mLk6ujsr9oeN7lM9THjNrAKqm54SJL7WBm0
Wy3zQ9bsy70XHj0bRN3/IBMfZNhNw5cIA5DU6g/cb01CJEuOiN7d9NIVbYwrAIgARcKIV5nLf5lQ
cEMogwJrfJig4f0XdznMrZMmPuRB1886PyGheO3hcBLKXELiSpbJDtWxaXnvxpfAoiBcPRS3uLHb
rzdmKvFCN4sS20FmJy9++6zP6EnSJ6AY5WYyPIGWjVtcv9hK4jJiDMHEs5t7toEIPRgVaZ/Mh5FE
M4vFLhLRGLgcVVBwKOimiB5rY6i4NnU2FixVs/jftClkgKfnKhRHRcNlD1stlASUcFYEI3oUikE0
nMIE/Ra+fz2xWP2WHXzeQyTtFssVqsiEEOJPcri2VpGWyRRufQJm4q4vcFGTHguEBbJYatqG0ZMs
rrRIhV2QGY8UqutI1CGhftYGywLxJbJsWQLOUcI45TFCfz9u7bbBVr4qzr7iZmFW5iULVvdrKbft
OdBLMCP/0tKC09yuWmENUwMIEtK7gIMJPyAtWAuJBvERRzzgvpN3tfI2vj8FEODDPcGrl0IwphCg
l+Adqs+bOUFj6+PxBZEbTn4giNbxpub3lNJSHwpunUQBbwEukPE/5fb14vetMWQHEYsoz3WJ9MeS
RTDpvHVGVvjb8AHi+Pu7NNOu89DRIUtjkTkBtB2zd0X55fxSibeOhFNukBWBOe5CmGTQDMsM1iPv
X4eYoSQzUuuK2e7zOvnQu5+ld2kUH5m8+XtS401teI9hjuYFpEtwiGXI3Nja8IkJkvRSdoDIsiRV
o4UbJRfU8x7l3W5YIyo7ElBPfhJf5upR4cRcLAkfTVBnlflanaxXL5Yg0O1MrzDGkpZV97ry/lXw
8svWBqk3tSD/krj2gvR7TZchkNZ+HArUY1Dl0oP5Z3LyckbIR+fW8wqDOmgkyzGTN/0WCdmdkxEw
69jmg5x5wCQYjTeNQAxv2ZMkEvxGxWHYYpk8eQTFQkYLfUOmGkFzYBMrUA6DRa1TJdVJ6gxAaoDT
mL5Xwaznn1ZtPzyXuHaOEbTE8QVZQTR89ybo+AGjO8yLIJLTnV45OEZf9IOU4vnHhhCJY388sjM2
YUPfurfU2Ut1RO1dEzQ7OnICCLNXG3wJudzQINHeeNv7WMCWkr03E6K8g7zbOgA47vQ86rEJdFiU
4wCJTVerQR/rbjbtKDo80hoIJnlqyvPGh/6c8oyLZrLnuXvqBi5oiACHmKy8frmqGeBOxwe9aSjS
MSb94BCoqMGh11vTlOIhGJLsuLbpw8LPEhBfw2Ien9uaZ73YHwdwZGe8tEpUWxtOnT4EVS1mjnWC
ed9n7VUvepieReNlOgyB4o7hbRx6fv1LYk1KJHx2mYTe/nreURgDC8+eClT0UHgGJSRsizIVsUwA
yiOyIZwdWpusZ0+dupw8TZ0amMlDt1/zQg0EmyLrqI935ElvC0y1hKJB45N8g9uEWtLyhpKdizI1
JkVd6Sgy0MdL9B2lly1qs8yz1os+tYSS1qdXiNqG+Qld7HaFVBwSD2dFbBsy2JP1nDhMwK2X4xHy
9VBBUEi89jOe3hdVyXthhHqSpKYdqakPWQC/K0GrmmB0aHnzRNM9JYUgxa4v7zBucuKpXl35izYM
MlsE8TYIo7Cs9qmUIbSDrWnIa6iO6Syhf8Z3xKvDJVlZX1pSfdWJ+Gp5Hrb0JcbKaSXawuJE80uL
J2lyMuFnJzUYguCFXhUPuJM/HIsmJ1cHjv0n5+Mgu9DqeU/z6UICpb3kXpB2IzNZDmQnPcDCNAVZ
baTw0a7dl1jfXB63tIcHVwseM5yIex3H/sxgyPhv9d/FDwG/8K2ryAolsZ99luGVKqDljnLUc/FN
53H+OYZga6WvU2JlvSkQuKe3o/MOeVjMq5C77aIv3ssP/FDgs0wSbkF/sgl4nro1jwH+pAXZ2d7s
MTASgVFJWBQBvtEdCGwzA09mBRC5WcyoevajP0UlZl4t247GYnb4QvzX3S7gYX5ePwMPD8QZWih7
qH/djWLR4Z38ZExv3m9c9CfOUrHsbIzICV73VS9+9PTpkHTKAmfKz3ddCaZ1vLkrfYYcpDP4Dv3I
JQbkxi2PvwFGwQWn9HwghODZ5v/gkQgFo+sduMYOzPsclrq2mJDOE7nCpv1tjefbK0q62RkfUmLj
1yWeOKFecXfLiSCsDPKbAH0+bfIOdTZQkOBPgnX7g+Rix+MwdOoK87Bhg6OkMPdifBYgoYonnU9h
dbzjdT6KQU4G+USkgQ62EiWDp4EHtycXU0YN0iL1uxbf+WubxVqxmZMhKXZWTwor5lKT4B/GPj+8
ZryctZE6BZN7FE7K2r8IlvVwsl40i2voGprBL0lw2RFVBu9ZjTjvKVhJ7LCrY0+uXxpGDtzA9USM
8WcJZrh1+nnov1V0NX3v4rP+6d/Bm1yRgMZXu7Jh20yVWIShGq8PjRyEVzfRpnv2OZGQJeyRT0jO
Efn3zDOuNYKbwJfYJBtyzLZvZXmMM7by8XLDe/lMBnt5Kf/CQDHYpAlp5v4An7qlAZAElgI8KVzu
gbSJO3XgUT8LC2b96dyn56EfKZJRdwRpGIVEnfU3wUTs6gbx2qe3wd+AH4wrgUOurKCdemTvzYDx
cwb+1vwaFfQKUslwI8m/hF9sF3XeRsgGoJERZyjrAenQWLr6HSFHb04fY9Qa8dx+U+wyac9VWj4A
scoILDWS1SuI+naRis4v42TVGUkCYsA1T9bnCnnnlEgeehbJeVqdN3px7CbzyLA7q0Dha/TH1i/Q
N80Qxb7kjaPTtPCzMVVmURPoIV5ThZZjzT5jQf8geNN9mwfupeb3Co6aYDwmeDKYPSXxnMKf7FT+
+JBMskrWRFNJ/GJLFDEUrEc4cnIkSoh/I0yBqHUZ6xP2haRwKA4NS7gMQVCL6l6NZfM5C3mqg6SP
noDMJ5VM/prHp5ZyP5NzGq3CgXBdxVN/RkGpGYWZG53lxynconYXJz0mjSVWHgmqlSzUvizfr7By
CS06UmRox1Thj0lP/Dm4p5Fx1ahyA88exDDTXYDyEb0FhS+KwWuLBSD8JIR+FQnqb90YAOHynL/t
/s9XIJB1uWiRV7pjfPgytgrySriHU980497l+ePhLZn6kRZ7i88fCxXHFBB42LTZNBJorGhbwBdl
V5c50QwhtUrJtlR92YtTmFBo6+qTlEaeeBYhJAGTPHKzwe4sVbL9iw6Q5C90mWaRJopfx8GxYStP
zomMxPRuzLWaVSQPgpvIDLQcaPHo+JX8InG2VuGG0QqE0tckxRZpK4IKOYY5e66TKMCoMigdChBI
s9A8G/hzB3c4jTrLlyJC0SoUTPU9+S5asbn/wmnKXD6T2nCOeyOi3TsA0pZx2qt9SACEC0x7xagC
bR/0XmYKk7tA6HOp5JiwLj4Ezew+Inw4J8RRloQIO1CPI0os+A4Zy1gDuh8zhebfjqB/ckjM2HwN
uYmvJhfRLHTgIvoWj20LCM1+C6YnS3PwoLmobLCznIsUSwtUuY5+GhvgogEexjVxjE6zEObfvshz
GyuxizgA/0zB6m1YC9ONNWQrVQyxSbJgNLQ3wigWOXH9migvXmFK7+UC8SprlL/J1zjCCVlXX8Uj
lldiuvAQXd9Gw9nxS0rJlITsrs10euT8ipB11EoXule5gGEodadJRiBOoRPbqvdzTO+Vbpi5ZsHf
LucPPNfwTVJcIL2/hiy9cUKgKRoX/713VUaEekkv33t9/l3xOpGeppa5CJmknJuA+KtzUMCDzxRM
p7JZ4Sh8gcgCSb9OQZmQgutt2XO76E+lzEaxfNHsr7LaI50Qo5m0e/Sejq8o6bCoZaZHhqs7mie7
GVxvMQjVQ1ksvKPD/LL9oXAyZPD2k+3EyIvkNRKBTlhmP5Muuj51LekddZcMktO6srsms13Z7I7f
n6/s1jWM0pkIEvknJtUdBXbwzvvVNl1PsOsOmchBPk3hvom9aDI1oDWVdWTc0tIosdwchhfF94F4
3Sdblzl7+CXM6U/bqa5qdgNzHFU48s1Hlp7BSKw3hI/VZ7dSd/2X6mRSWH+kSORUrU/Ulp+cgKqc
wNd5Xus71oPOggeI5lxecqyZMz6Abt9O2GPBu5pN+G/d+H8j3XUvkbObtpW6zjV14na44VWha54Y
3OnP3wvSs0tN4knAH9R9zk8JN0sbIZqR3z/5LGsIh8ICs8ABJ297N6Sh0SrNKN1yIwGVF2xFdfoo
6IrAB5Jlv6AOwEqq7K5iumaYC6tOm2vqEnz1tguN+Q8BmV/8wcCHmZ1p9dpVDIV3ieSZDr9JohNC
8A8ZYEO3BykWi1tmBATf1d7BgjtY+jAYCLLepu8gB5vhOiohln873mFkoKE8LY8rs79yRx+R0EDE
6aU4YREqd+Pk3y5/SO0k+EEnGzz5IEmULwZEk3us9mpV79cvNmBjeP/HOYi8P6buxjcz4xA13f6g
ztchadFqnWYbWhnb1GKwiPYXKa+ek0afNev/jKt5zp/jem//spdxPqbws2I/WgGvtW77beq7BK1s
ASyCu1JIFh1rQXxQiunfDRIYE2jua9laUSeyXmFp1otyOinxa0PmRoFSrj3P2AS82JI0zswHrMq/
pZmXjWibPpnZGCYrfuwf8RQbRM//0ZkFobxiQ8vzMAzb5LFOtC8R1G58ssh8NFQkFqrDFBApLMPN
lVI1fWsLpymZBiETthmDNfuBqu3SThJ+r1Nui+mjvDvOFyCxyJFq6ES+YSy173BAbOy3vLWavAgz
jUkuJMjZlWi03dw2ZReOLVBpCR4SxbUGMDdH+54RdDA5cOOQpJChNqZnLgxevQ2NcMCicoJ9LZwJ
8RFiNbHfkbOUBGzMqbc9F/E6sXxUpf1ArfVx2GsOgBlGwVIC0gsby/4XM2h88dHgM4ukRzsYde2T
CfAFvJgfIBUZe6kSTULSzo9SXpunbAUVFCaQCqHVDmLfGVcTqHqz/XFIEezDCIZAEg4tOaranNuJ
bctiP4rmpq3erdKMi902VrcmpqiPC9ClgqfHPnD0pOYFI19E4lg2JgB0kgMUqtHzNnsum1iHZB6q
g64AvCcyZ1hUBsLwcEbOX6S3iFa23dx5hDNBvBdwcZeR7c9N63et75Sd7cTcIqaL2AUf+ejq3eyi
kt5bp1CZl027wQN7XeTcvOlVwWehtK2OyNIc/8lkKzi1fHaThHskg/gobf4jZj9q6EC/MTn7jQeJ
aV2MkRgCd3ybRw5FMfDvM4NNJmMhCrmw6mnPhLXLFjp0NrC91b1J87jgVJHrRu0coDUedyNqQ+XB
GAREF1n5uDApLjLUwjspDpLoKf8mRlihI7/3sxwTopBjdEimTqrhvG25p/GvsZm0SgL8Yj5ksG2b
LfKx0/7cmrDdPbYMV1JY6Q9A5CKf2TdUmsEceyCdtJklOAkaP9UMKCy4usYdQNjl/Rf6PZ3jVwO0
dRVpOQs8iasS/94wy/5+HabuE6DATarZJlLOv5wUQz1RAnWAJC1jihDowfIoZxgwRIlCQxm2DMpr
ZbjXLH/ZlwCu6HsOARhSjlGT7gC/6fQ/DFiF4cv8UdflZx6H3dKv+XZc/hsgZpJFbtmGQmFdOFTt
glgrUWjFDA2KDwhbfQotRWBfAMR3sgO7bJciKKz0wF7/gAfo9hJMSSkvrUVaB9V/5F+Oih7avZEC
KpQR58jNm7wpooKk3FN1HXQfJdJlP+VzwPBj8bEoaoDXj1ktxojsx3UsGwgsOkt88JWmdt4mcEtG
+8AtqC0rXDwBBbibsYgQhCOg+nnkqnASQG7kFr3RItQabc0IuejrHOQ75fM9yeHBa64ertcqdcUV
MlnmT+6e+oXm1ZTc2AZzu32G2H3yluiPvLM8v6MRDiZvHLj7EsTrB/gLEx66AXpaWIGKeFWn7LOp
cKsXZMqk+vQiESU+dzixzEjEJt+GuqBUJKh7+dQDfem9Z9UnEUwTTNKvirPrqqWeybgyO6hVgD4L
Pp3aXEo1eRfE9a82UVnxEkH9/4Xsh7Kz0R557ZrNJsTm4csk70P2x2/28YFCdcV/b1O3tT9SDErt
JPPMtCJikjyPFDYPisBH9jTRdGg9cNSi8F2z+2J8ZT29cUAsUXZ3aljRkFJF50j8T6IySXv9e/PF
PnFWhTGkYc/RfVfXokeG6XdN0PeGmgV05qVPWe3ZqGhTk3bKQwtYy/lI63pmX9Q6rA6q0xMrnrLO
QrqJtInEwSDZ5hGZqqMC2umS2mHJtD4gvI4lC4PlYBH1mT2gA9Qp1cB7QeXiA4ju38lCcuN+tgoH
2xf/cr/0ZyEILAIzgGU3M0vZxiL08D2c8u2VnVd5Mw2Y0xU2W3VwWqc9eqnzEnbksZMmjk+hBxcf
qzUlwxn3lYPURNCVh+niExajJtcLxC2q37c8oHx9Z5IeP1RF/hYoCM/CoKyw/rqsAy9dNqmCMyH+
lMOw8J+w1BFPn0lQiTN14bBzeBKNqiHXVo4CtKEixNvr3+vbmVcC25dOGImYU8Qd9JKI+NPr1esy
tDqBpKQ5I16OBq+7eB7Slhx3lHFDPZgVrMkpY3Isiq8OKi8brb1/Bc/J3FUjx97Q8XEwoGYiTg8y
9NbMpgZkHeuo/gDta/J8kwar/x8KqHx6sYtpLXpoDzRTGApmYcGufQrya+K4mnXJ5H0j/9qSopcr
LGDBP0VRLwsJxAxKy0JUFsXPG2T752mHYjoedqaPpytZcmOc7LMJRjdd8YntdYIjlxt+DwQjXaCF
2ZLp9bpVSoQV55M5dZ7ok1iBKKHI2QgYbGsz/Uyoh6ehANydP9z0H7ubd1jRLC7m2rvnlSN/EgCk
VICQVEJqJzON6htDF53pDFOAUAJ2jBODQpf1J/5rS8RsON3rCqSk4V4zJ9sWRoKJm+cgEWwBlmVZ
VBAMNzGZ2rA+9uTVP9ExsRDo5e91IhTgUnZgz1Uc5U2y9rr1Cr1cteti++ntL4vfwpR68Tr7fRCw
Mv+dJHIojylqxT2g662w1J/b4SxSN2Za+AyON17GcJV2B/ZTWEtUMvdJwlChlQuzffGLWz7MNCtl
J9mDMvW3+SxMd1Xd0Jyz7lnSHOVU2QPxFViZcDlFX4dyu/X4yA9ljps53ivTL8YX42BCaegwIhII
PbtDzTU/H5HHqcBjitLEz//8F/WiYL1pmnbKwgXI4kNLE+T+BifHUtmOasJ24E/xndmrzEpNR9l4
CznBOqu9DnQS3EbqgBh+wsWbJ1kiLkDRbaTSyfDYDLo4nWjjVhJxhSr2B3MQzp4uekj7my0Qc45y
2N2sxm85zY9hzvFEG55mZ5MD70bfUz4ju4/0eq0nt23dLZbjHnokRY3i00/z5aLGBiQ8y9n1NDq9
zsQhs5eZ3/4E1PjMXf4KYYdDAXwCgdLdVRoOaO3cV3gxaM+ucwFqVhZrvpOeOuSa9KYkrBGiw6XX
mvuuWQbbkmBhwQMH5Qn7P+DTwQpGxTtJb/ZxNI0Ifyqiw9f/Q5DAghF7duo5oloLTUE1TDczEG7D
EtYucLKGgdUOvZRqCZiFv1U1pWRGV4WCgxpwGBCkq9q/WiLyqW+r9TMSupDf1+hv2YmGu6u7pOoq
4lZSy3630rVvyJ5V3EiUt0VKgNYKwXtHGLTFZSk69sudp5ck/icvvf3X9QuJJrdUFdMRO0kYzs0L
cDtpolP/7oh/0voZqYBHwpBWcJ79IEPI28uhEXtu+obVfwiXuQHGLk/v403Q3esVR27KG50Qosx/
xFlT6zsJl/jumxbt6FktPcwCrjYm0fNixSS3F83E2ZdntNki/JUWHLyrKubvyRcobUM7ebfiFzru
FB6MTSA+/mBEMTRfKTdkklTXUvMemi13fnYrxFRKuf4ikzNsP+Wo9avuz6ZxeHc8uWHuvmWArAqS
KEm2/5k/F61f3IcnwESOhGDBFzvKns5LYP1gaKeWAozLrfKvNqdShJZ5oPrwINjGf/KxzR82su+u
Z+4ZLGeT0JbyvVik5zZneFWKZ40/eJVp+PAkWIa+0srB7YE2lLTxcRogHpt9qCKlq/UuqKezG6/M
0Aij8NZ1e9d29MU1nNrlowDl1L1VeeohEvbJrlR4Gjph74HC6vvnE0xHD7V2lNaJBflT30lrZPCR
YHh6he+Z3Am7DLv4Y+Fsij/cnQltG3U/zNxoaCgZ4AEsRBt6QopzUOHQvVu0TsMxkgxSoNqxqJqj
BW4erLFn5Rz0I4gSvaIbXnFwKRS1xlZa41I2/mS7ckGG+nE+J99i9SSW7i/As+qKc/QNnOhRSk82
zs0LWTzUA04JFhve+GM20VKnqyGnw6SPu7Sg4143vVu93XyJXV1SVtgy9E23lrO4sikpQzAAb/gU
QBqf1SH8DkKyS7mgsqn9g7I0ZjVq+a0GO8n72CBorB1pXTpm0idG2418f06Q1XZ7G3vFj2FJ4Ti5
7c6+wCYWGNE5Scb0PWcmWsgU28WXavOWowEanmndgTem2AI+oKIHYYN8L4jItYQZVLrv+CfJF7cV
0eLdUZyeCzXDI3qRpRLO6Uq9SFhGSIM5M2HH0lTDgpm5rVZYb3TmIr7eQIh8RKBNQL3/XjCs1RHi
6CgedJrSvMikgM+aKdMtDFaehCYguF6XYgPdOLTR4VQAhG6SCmuA96oKT/TuuCip6LA1xdyBxMR+
DpLhijUI0Tv74vgczkYywb0G9bzYFqvrgKh1MHdD2y70bYYWzM36rPFJJEGNblv3IN4mn12akAx9
WSDmAb60holKsv1iXZiNSVm5CMnMwOM92srslXOMYCZSocrmfbgE3DS39rZCI40GUmsBbEHbKQZc
IBiva6mMkesbJ2uSZFUMGYhoLI5spolCdCwYJLzt2FmqCf3RxHjvtb19CO6y+ug5mnxYTxIMQNfk
3UVLeyLTCryc3Uoa6VRUI5Okxn1h01+2XUjXsSB6/VVeooWwWEHeCDs5ERhSEDUmmuVjHb/oZlV8
LTboZRZRiOLh9eeGWgJE+BwMiW28ezYPJWKJ3hwRINWFZCNcB2HNiW8hTLQg2kxrKu7GMpQG/K+c
Zi/uG3epkWwF5CEmR9//MnuHuTwwxqdD/kLR9cmKphthcNvjqVbGpdIDOuuZSNct06SXnmb8tD99
L93SgklzRi1u5ZQIKV01qdU1OxaImKLTD2UxmES+IPAK1iRzt996l9TZwWZD9MEZ5N3iVlxy2tYe
bZA5zhUtTcoGxBDvLKcH0oC2TbcChEXtk6+xGvViFs2zWh5PHqc0egz2/JZmU/6kZaSqyC/l8Pqe
LJsTq/+M5BiwaP+ROZzNBkDOq8t3/0Xkq5W2CNDCQJi60X92ihXprPTlCzACGWeFu5q6WzfPtH0Q
zAcqITvbedQK5NlNx/qybxg9f/vkufXVTshnNcBxxW1SuU/0kY4/2H+iDUz3+prP4YY07Lx4m82j
BLbd9+9qknekVV7ybp2jWbEA0Xxzfnrs+Rp/N3QjurM1yWq1z03fyGTUbZWUhTMMpKJ9NcKmi/cv
/YUsdA/SYFUdsYtAFPNHYYy+/dd/sr+/RyIkhpzcbwSZOeaBqu3zk5d0uZqfPsWzic6CM8ImCdnM
ofb+gL1anrzGcDfOKutIlo4IiN3vXcR0UZlPCid5SopGpJS8jJAlUJZCNatF/WCvCiIpcNCekFGg
7j/tI37PLpxIfXlo51/Lrck+l5YKe9ohMRvp8E/vr+jFeWXuWb+ShhiiOnxF3HOI6pvA3447Ypjx
4PL4eQ2AG30ueJ651/Qs0FxhX/KYXcMdNhPEhJiw8JhM1X5TKxWKe8NBXS5zny35vVvOCurfJMJ8
3eSvAFghii+wGoZJtJlfrQNRod099aHYasOxkt0Sx70IeuYJp974nak7aEmr250MNzX7zFtFxYjv
LoULovY8FxGpTbFfQiIVvXc3Efv0Q1vabOpr5WYnhCU53Ux1xGdIvm7rD3WHDy8CE1PIvWWUQUD1
of7d3akRqDjkURznyJ4hdLlcMRO704giCZBgSEXh7V9kOPE6c+HtKIrSUi0x6rEGH6BufmK+I34M
Za1a7V0sfUg/tGuU6YxRKJhaWquHFBo59wme5aKo/mpzRoThbsvY+gZU2pqFGmRaVy65vnMGwmmf
oPoaceCEMVu0deVagtgJcbFBwSZyWiC2hRbO7erwMBnLNoklhqzsHXXsbZ+cJirntng8zqIDaeZH
tXVE8mlR/3AaBc9FFAj2iO1TuZ6vYnjleZ7rQMnMMJCtqCW/MmPSNuUR67BxSmkM3v5OXJBe6gmB
V/iHFiD+kVw5rg9MESyAr0SFYAc1q5j3vkjdWtCGKNdPdnC6RYE8KN9TMmy7nZB9+rQK6MkogB8l
j5rNK9N7+8WBLCKlmKSy/TnEgn2JzTOWeqrO3MONwGtOZJ4F1rStiZMlMDLj1T9mS2jl4pPjClzs
ebprJhXCR8AONPwJCHZGbZe/4f/79FoJfs2f3L45RTqE59m2Q7KBd9HlANOPnW1yhGZmjHwPJ2Lx
21H1SfvsoSeUNaQFoMTD2s65ZJUGhuf8WPdLa8G/D7Yie44h0PTY2S5GiX7NF1chodqiCSpcp1kI
lmIZSx+G7JueQOzta4fMXoeE104Tp9pkchGV5gd5iNNFVZLSH/gs85hcjtsGrYEK9tVwdO6wM+IP
/bAUaOVQe2fXWK8k+uSgXSWqMWwvOhZFysi5/M+eeMtPIjRFXf87LWkHYvPbS0EAfgQuvBfn2w1B
olxZi9MMpdcry4BDC7GAq88IVZPahDA7WUTVJgLKFFRPuNb4IOSLDsutdAeTmDfvZ2D51HDGzgfo
Gwm28y/+qmAluWcu4k846PYjGG9C+2PNJdtUu41HqY2PS14SveEWBzjEFabwJovViNlGxP3kygZd
p41d2eoPTtBocP+9NBt5Yxb+g3rs/mfNwa8vmZYLlRuQxDkvB9CyvygZDPkMHIpp18jT/s4K9fYZ
9Epfa/5R+cKYX6ZSqfEpNKKrMh3FIEdaomejYLfILmCGgxYdKsF5RKR62cDyqmB+uqwQdOyqJ46x
5VwuD+HQGSM8+pVE1Qgtes7vfqkPwI92+c6YIpFb2J1FK6TsOwGOuvPcyxlSMy2ar4LQb6as2Uxr
hRibI2Undhm7CyM1bNsEiTcOxe+lItVcLCvTioCTr7ttg9OAbG55ihHMG8S/8tp7iCiiLtSqMy0O
93d69X+LW7bv0vt+YJDy6VaixJAE1C3OtDIXDNIRlXIrgvymw3hVN0WVO69EkiMrbdQfMHDFF3iF
UsM6yL+qULasKtzHfbhCe3GB6zrGRJYdQ+mFAFKxegl6F67bgdNlPwPPeg6mbxavShQkyYt8Kzjo
qJOLoaQsmgIRLDyudhctMLeZYshZghIjyFwVjLaOtOO/QUj78024WuiaUY2AYBGhuzyXqvcG5Nvh
ehen22rYMavsICkB09LGQ5DWwBfVgsGX3rcQtu5nTjG0B6RN4NAEwm3WPQnpo3WKzk+jZQqCzwHK
0yQvXWGHDrrrd4r3SR+U2gjz2SIkHX211dDCH61fy1dXQUVge4/712G3tkge671+4ioJzPrzzljd
dtzGVwwF6y41nkSvpDnrtaDfxHwR5eeO1d5+Fn5GtxAdEDdYkWebu+O7+gwf6JCkpFcObW29+V8e
hMl1ryHB00q+xpK/YLc2yhujXQRgqWMQt7z3BSdQhVoWsfojhC4FoAvIoSVqbG/qM/9VwX003Xh6
PvEKwVmLv1/UH/F+lFdP7TXQErodJQuZGad4SG4plrtsgUNThbDJiDZnEtK2wELuYV20jFzqm98c
OavBjB6E3lmE++dXX9+MWvc6K1PnKsZtV/k6CKzq3bl1T3681jV57e4XWnFzXh/h2K7y7Eg6fTjY
dmsOW6/4S7511iwIoc8LGqYVLcQWY5PrRm8yGvMamsiu2hYgEc7azZZkOAK8V5lmL0DYxkE/57zb
VBV3fgYx3wb7TNv9zBwQyN9lTLeOfG80GHqnOGvjDb+quf/x9gyn9i+BpRojSfbK2reFd81Gwa+T
Pt3+ajg6tsIGHTXeWbFh4OiOe6MnmI7G3tZJKdWlPhoz0IhYIwnk1mM9OjZLWd8JFxAbJL3o2+/u
9UadOiGkLxelY4TB5t8ReNElVX76J/+JVkP59KRhQwCaC4HhE1If0xO/CiWwpORmF2uoRkdA5QSS
zcxbTMOQN14sNHrHTuBg9UkP8ulIfqrecGrTTwJF94sgwlvA+B2HePN04llnqqkdnPa7hgSrdkgs
Uec6j/gFSi8djQk8EUdPwrnpYhyB4Yf0esUuYPOPE8PcGFP70o1UV1nL6tIFiHQf2GkNdX5SSDqE
vlxDVqn2vm2W/NS1V9YD91lxuGblJ6dBZ1pREwNl8b38irq4kodD1DqWN57PNqxsGr33UmP6Iz1E
c0+n1l1EzmxtPLRKP/+pHg6+FBYRa+z94vpztlWSZp0RKSjw/fkCwJynflF2KGnK5EOmXaLWxrJZ
x0o2Cv6/Naram+EPzGFnFHO1ZHuxssVAsqQQ9Q6BVeLtplAoCL6XeJz3dqZDkm5s55JveyIzuF/Y
dYihlACqUX7UtjlmX2vJ2DXP8mPhILVfeEfDGrwOaXuF7YqMXNZeNfNGJ9TzKZaUuAyP8tes7efI
YofNp3v2MLUCAHOMm2bbE94HaNJAgF06ElWqwMWRrrZb/2rSG7SF9EjildE6OsZQFB9wMdLNyy/l
YRW5BiIH5OSsFKuq28qEec1fFhB51JGf6xNX1Dx6sRrC6vFjj6mEp7f6IBVn6g6pXCpYnrn2o0uO
Im9SDYsBpCUKAHOftQhEKbVUynBYA5K7llDlDaOkpEGXc5f2FTafgMMOIyzbnT4ijtIw7K+gW5v5
/xh2HkHLrCQ9lhLY/NnylSSqsulS4ImwyKNOJmecXPt2+0GVNv1PxZNdeJxDaOjSEdcUYEb/RYNz
2Shcx++XrM2jwG0/qqu6X64Dqn8Hh9tii8GF+WU5USrQNGX7Ox5BubGStZ6xEj/sSk9Up3lWHKGU
FGcx51xh6ue4QFbaFFVZ8rzl74Rf4mu1WlLV2EymCi9v87P0wD3E3/SJ2C4wcmlQ8FGQKBqEYQov
SPKDWK2hC/1yDQ+/os7013aAnj8o/j7DCSZvrkMYM9Z1UyChx8/3UsI2Fs154rHWEkbxhVKIcz12
hBbrPqVMssCAz7hIik56szAxig3WHaLSitDkZDTNoIGPzgl15WdcqYH/TzIIYjpS9OiX4d3v3ykD
1gf8KmpwWmD2JxI457L5+lxW6J+60lO6PKj1xIDFNncf4NLog0c2xWqVci6OGI7CmbCzH+ylZRyH
8RSmYjwh841TNZx8LImymaF3d50k7CdOXYtn/SfVwcVe5Q/k0AnDL/404pWiAW9jzhVMCn4V5e8t
7fDtJB/981oBfWzlHlRI8gi9c3QSbqv/qDGyuhgv4i9Z/CHG+irhoLwCaoKkLhqj5KPhq+WV5s47
FFAvEomq+c5cLAlDvzp0Qlt+IF/cTAKZnA5KPQb0ngylBlFN76IAKAw/ZLOi+0NbB2DuMTb+WgYE
qU2v4k3eWsMp3YN8Sqymd9qiLghsHNe6iAEw7DnxoqITX6ID8/6e7qvsmYk9gHFlsbMybOz7/k6L
26Sg5+erb4idzTUUvLbKHVjXOICsGH7HVFH7KQJMYlZATjThpIr7c459Yb+cw+SvYeuvlI9L/lC1
6h1CRz0k5Zaan8Jz6Mr7rzr7mnyqcUnJtd4BoehprL16Sn0g05nF+25Dufs5EnV0KZfLURweGUFM
9i/kwdUUENQm33+ZrJ6qQbl+NdwGpJqe8o8ftZTVs6euoVmTZqwOCkSRzbnA2PF3tHQ93JkXgJgz
Li1NGKBHIGXqXBKpKYY9HyEzny53vKVJdaHko3B8WRpGH7Fja+Pjk10EmeudCURRjSpM2TsTBbGw
A9zROABHIExRGWSxRQhsTR7BUA3ZddCtrLoEQgnKb3VVWytZ8KFhEjBVtKTA/xgqiNXO8T5zl8xk
wL8Cc+sR9dQcfzgWlfUxeOIKh3ffjuZ9EMH+mbp5Nd/TMofT44BulW3T10DleNW2oHMByFcKKI+z
7k3pPHhoQA0dZGsj1vWKsEBrQrXaoO4t8PHjCRhGSoc2s21upQf45j8CeVuCT+6fAe+g2AtfUlTX
s6u+VdMDcX7xh+0F9zROCNFU6kW7uZdD7V6q+28gIr3Qv69p4e6WcJOlFbBg3eoMvFAzSQ/Bt/fL
8YvUp3u9qmiccJYxPhr0jOR1xYOOEHcqpPvn1ber2qv65TTwpbMG2QQ7FkVY+TXrTUiPs40zsXeh
qmeKnifTZ65oUnRwoWxMesULMRCOA4/bgvXNxMvB3s71HcLz741HZlMQX0BrNvkx6JcyhrdKXeP2
sGydxrVfCAZXDX36B5RXRT1XoLuwnjkwSAhEWgtvSr39tdmoAgxqvyynqwuLbJrBLQ9o/DUyyCSF
0zBhZxBoUghlSKPep6exOTG3nWBJvy8+n7sXdV/yizAPy6RL4jNT0Oia5r9k4p02DiSH8wL+ML0y
dwOPGO3Zi4kv9xxToi0yW5KXlrPemzFKh99KNFr+FK6HETyHUCKA9XVefQq7RPm2ydY/PBlWAHaY
U32lF605zssKbhUJsziXhS3jpO4sSODKGcrGrApQy3dy8GdPEPvl7xDlDhfPiqWJGXI9ohAwhvdt
BoIiFnspKqJUKh95+cgJJ+KO6sd4VxrDod9fHqVmWXH0cTTosi7NN4pZzMuCuaoO6XAGCZLE/LNc
0zzGH+feumy0UuhEho/SFHiBNbvq9sPKhTSGdrX6nWrp6DB+C6I504y12tJiOqqA7585gcahzPo8
XJUkOedWHBAFDgNMOsL/OQRdsdA4x/V5u59Iz68nbEe8H+UAg9EM4v6jRny8XXqplDIbtSfFqVxg
4QSDHAVKVBoW6U5+ntBdMDzBVCrBTl90JSJM9RqFRI734tng8kB+3XBXferD35Jvb0fVAKWmcacN
CvUWTRtK+1FDEZc5Rkl2AMrBjQCscvgRfW52z5dgVScm0ntFWMYqf9YLMBcXBvgsfwypsD5KTJXm
XMZ7mxQI7nNi8LQNiEqBxiLRu4xmLLvoz9mprL/4sbVBoheC+p1OHnFRQ2+S1JJAuGMvHdsfMjmn
3S8M4jy9DVIDa0JbBkSMOwnItUovvBMBapuNPdnre85YdtDtH/JSGlJlF2gCTB1lB3QNIKlw8z+1
yuMWnLydf0oI+HmuhkTtk16aJO6lzzsMfR7H0nlqzmWz1YWd5nm1M+tlO4e1rBEFp/G+5PpQSkOh
ZJZ4ZVzW7VRCRTIwa4d+36sQLrJrO+ISmBhzLHvO/GfQTV3QnPnLpY8BVymE4OcI93KEZCGylDHe
t0wtd7gdAEwEOrW7AKY9nwHHrLxzgpHLlBVGNuFZAIP8G3Q1RPAjTBcb/5kijb2Jh33WQgSh4P8M
s+Krx8+fqD2I7uVHlRrmPkESIGTzgplcaLUP0F5K4s6KqQW4jg9BAE6/UXuMZ1cdR5D8mDagQxmT
oz0SHe0LQLTP21pi27LLA9NlcdDv5P9utbxgNo2Rt91SrrNOJnUn6Dmzdy6MDvBL+EMLcxEw2VFM
9OkqeOPMB1EX8QFrqASxOEpzh9brcPcoPUB35OpwLjdahbp06Z6mQPCGJenMhZ+DVZl9qrXHu41h
veSxowpCeuWT1uNq8vDU38juFDXTqGDWockCaQZ3bkrBT8OANCKfWPe1oNkkWOIXgtwLY6Jp9bw2
/G4vyp6c5j+exMTmquvnQR6Jk2JJsjJTDlE5sJ2zBnfM3Zn9++mNPv5G73MJIn3+rmH+JOYu36w2
cmfqXBpBkh0m0tJnIAnRpuu+ycRMp0oR+spH3NvTxJXZuJx6mF8WXa8y0wJe3Kw1uaXGmlhWp1pO
qW8Ml3Rh/yuwMYtBLWa5gs8/ai0QplF33nzPJbzZKpTeyQCdc7pHjyl7A4B/DA8oWrZ8Rcoz8In2
6SmjpTrA4jRyA9eMbMxPqW718VGYTi66F/TZq9lpJaI8nJIu7tqy5Rf9xt52y/Uf49UloALJHUMW
cZoHgtRJN2TQMGeJG1wpDWe4fqMJootjYAGnGJ2rr8sVzTFtLoql9CcMEBp+I9klYUi+geqiIAyE
tj4PWui4AfCCwSJP3Dl5ZEWmEiUmus1gmxtI9e7aWYE6ENxXVMeoicd8fckpJf/iDg3JRZmlvdMK
GBqNTBg3jtgsit1ypESJ0Dty+2DAtJk0IMUM9XXnhNMNgGgiG1ggcoYv6IDa9KW19DBgGbjBZtue
optv8LuV4Ib1hKkU8POWSYyvlVvaPz4pyuvF8mWHuEC7j/cJ6cwyTkdIlzGgRbLM/+ZO4pLgYEj0
RHvVC0g1d+wlln1a6+fzGVLSC+v7KJmOiABVl211LAYZVPhpacfioR2h8DiEIUGefb+lsT0w8GzJ
HfRpNWW/wqr09oPo3pgBnyRtGRJqbxeU1OmGnUI8lU3Z1Q3iAe4asFkDil8McHux9Pg2X7m5qGbi
W/aGJei4m5NigwwnPS72HuVUoFTU49rjsD8c2M4UqmJtkkI6s6rxQ8r152DeaR9dg8FpsUWARysD
1yMGsGMQopL6WWcK+WEDw5DoNOS9TRekrN/XFxg8eX4XRvNewzunWvrrpOOlnGx4QUCyUHndD+x3
SqCRNW5TSzcdXlaZtCmhbTeLIAJz+N5kyvDKbHVuTwzZTvZPvXQm2Sx3TBfuI9MAX+StJ314FbTX
hgRCbbD7rSN6AE0eYNDbz03IWp7BtUJs2O9y5ppjUfIAyn78vkl5npUkH5j9K0ffCPZkvBYua0r0
G+1cGYQTRCO/KF9DSNdVNgyJrW+bTWHsbEwR8qYo2/8/yxDRcsPsUgNWh4aH6m3YKUR2NpZ+neob
gQMkUN2oMjtxiQITDcw8ayF5j2Z/lm+0vVl0/EppEIzd26+f6XaPB+6YqUGOkc9QylXo2FcCER/k
UZzffi3s5AbIHhr/Aye9xaTe+QtqPt7UfTdP/ikCOs1QGYWy02S6/9LG74IapDTvpchzGlvtYvPm
0Oi/DMu3u6jKq+YL2ls1O4A/vXEpv+zfZjwioy0xDVESqJceNZAJFCWan8EHGbYUP9RRZWfmla15
ZczkkhiSWKFN1zgo2CUwjVuyPabGlGBeTT7etdHDtG2sPp6U29UEM+xj3l1s7a7IxZkPjzzTwtNc
mnX00xnPCvD5u9/5jL53JTUoTTB2C/Oq4hdEjGMcgOI++MsRTR0dfvwvyQITcAdAgrpDtwrKm0/v
GVqLt3sI4LjWQeqKato8fb8OLnQ7O4I3wa3G20vGtMZ0n+BhOMa/6+jEtuAF3WMeXoofjPiqdrU4
nyNJEYn4kkdSqmIFE3V+yByE24uIvsEdZl+vjmmsuWkUjQ6HykQbGslGEKCpy7HrgP0szib8O7+1
86lD+57jv7lsBxBPy2Pl/Xfh4CDTDpdQRfnsJeTtMl4Vp5/fftzawq+tUe51+M30fRKkYrODcYdg
63kIC0RHeUyG5vTG7qrFBYYaeqBOwvXyGUwp6J9OU/9xZeBJLaBhRSMrTzb7kUFeyt/iWPhooyzz
RvETQKus9qGwRFPEGrectVHFvmIhiQC/cLws1aZtfuxBSL6vj50wQ4P4hLc0TnQGFdg5ow9xIMWE
KxAzJ/m8J7jkOivUdt/EA8c0ZKzVXLrIrKrPZtuxaprLVCZnLVcxDfEt4F6svKw+9f1W7tQTok93
xhERqiGdp/xMzUiSNrD2bY7qT7SUSjBk5f/zP+RL7+/nCIarTymkMsSW5kkZiUB77ilf5kRHTr5T
hRZOAH/h2PtIkiHXftIEeSoAgMaRdZ+OEH9jCgu3t6flNujj2e4n+4nhPArw7Dm+hTade4yLipbO
nGqqtYY8LvXc1pboXyDR21UeGZCI/4vOYvN4eCw2QBYmijD7BMCxCPTtZhG5uqZyhMxcJ2U2xjAT
cObEVRvHaZEnqZhl2AnP9ldYqtAxOstNc3Qb6KAXbfTGYfo7ZUHb5tgp+ZqQhtGmZaBzYnn9tcsg
pqmgKAyEBnYB9+WphNrzhch9r6bMC4QDJVQuhqv44GkyhgayH1SmcQxrW2fly3sbdIRCQW8slymk
w0WKPj+u6PZwxqlyzXo+35VweqLP6dJAdg2ybIVx+WNja+/LW1l5INmVmgKha3QLL29b0mAyjBIZ
AyTbk4af3zmc3+tUjagHAO9rkycab0EclP3yf7KRP/S9b9FauwsHjTpLQrENUgerZzw5zCTlwLie
pOfW7BXtMHcC6PilJF125OjuXxpDdQdVRCQln/5CaaFpd7w0kA3t7tAwL1I+sO2Xu6qmCl3pjDqT
pe4kmnFR22a84wy1ClrfwJPmdl70JLPaxnTEGKvkXNhH7GzGsiO6LHhoCzZRjlmY2ch7FQDXfgBa
pybsX4Cwh8DAwpJu2XVyiYVYxst6zScEeiSARSE7w4WYj2eHbsg1Mg0Jf889E5kxG6jQfLs8niVW
c2vKoBo3EuWQNzPofEW3JM9OCayNshi/bpa5U6Xyy1/CQVniicB0Ibb0/rXr1KpJwy9zGqviP/qz
irxb6yo3c1HKsvEKcmp6FO7kwhEKHHoJvGfyR0aPezjiY6N41fHqy45e2QOn36TgDJ73zfLEPRxi
ly/4/3nZazFMMZ5etEZ/CElyxSk1IVe+Ni/wkO7IQWJxmSBP3fZZL7zgaHorA6bkGdXlbGlHspXC
Hg90p2grvTqfb6MHqtvsAGS3BnQa2nQGzqp7Y3CQRySlXUI/jY7knuC1hwXPMuP3MEQ7hQcwUqlW
BZ0vJVDEphUfxJOW33f/7duZCiZsQ2tZlF7D+GPYrZpBr5RE6gXFsADPFPshGtXd686uYkso5+3m
1Efeur4bH2caotOgZm24b68p9dQ0obUJNYLyLBl+OXB9/SWpNs2Tm6oIe27f7nrwvE5mXM2N9YQq
tNkjZjiEuhkGdRVoVrXcrnlIH9vIQfnREYH3a8XH5S8cka4Q38ggMksopdGv1BpzpJvnnOy2Z707
Tiu8kR0XI84PALwYsxKOI/4ItsV3fbQd/bvaICL7+GPAUNj4exrxLzlvpRt0Wcl7BiwcSz7dTSFM
xJ4i46Z50JOQhSXT71hg98VvqFqN4DxUIs4CQ4RBXPS4XwSTXZXG4fpqAmTbhnbHXcOIwrquqit3
Mmd1gtDDap8DOrz3AcNcY1f5ip+sEiesSMXbkacXrHalB3dPYvO67RUbyV1I+bkb5XX8lJ8watDb
plL6nh1weNsnsUpeXaH1De4VWE0ubhTyTeKBaEsNHVUncy6E4r4JkSSj0KkVvivDViAHvUA3hjUm
XU8Q2vaq8AV+KicP2eprmPYD7fsdRUBzCLUVlPMVzy6Skff0iN1wOvZlaA/DuNXSZaPSsxyHjErB
Nqlc2DcpyunOeiZ6BcRN4jxgyfsFPXrKejOHDpeUBQ7R8Zi+uzpV2QGkRY0aIK7xSd2RvYI9ALxS
+o8un1qs3XayvsBUu2C6wEGXZGMMgG6zhch5O9NuRZB2tH/BGZtGxrRLz3RQh6EO7QDlYrpUDltS
3cR1xuv4A/K0FFONYnGlcrL+Or4vjnFHWrIUlqDu3MCZqS8wxbv46QEc2SX90lknathRUaE9iphd
U32ZeV54jxddLaxV4zwc4i9HqmbCGySr1EaIA9x0CBRSRJSZaGJeI3DxJ7SQEM3sDaJlFhHYPjA1
NBHX76Z6efisfs8QPgr7mSqlBQ06FJFbrtEEZXURqIEY4LBs2pnTFZHfaanAkxm6IPXPTknqFQ24
6XnpZf+xacApBzP8OPGXCbtH48+GFnBRn62diDE+YJI+NBAfaSBeH9Gb3F+3Wce7CJVqMUh2UWEG
c+0msfHExl4EDnEJ2OIdmPhQN/YhbGjemy365fniq6VaZRlwQnzISu0K7f27yWRDO+XlvHrfswdI
5rzeDtiD5+CTW8MEqvvLcFBN+zCI0xTtIQVaFDuKiiq8zMw15CFPfsAskqoJwOFPNsNOveMZOo8u
9Zw9JOeeZHxn4fYYJ0mGwApDEAHStG3MWZB6453EIFW72wuVDT5WweQtVn9QSKeKeSPI8GxH3T90
o6AKO8X7SetMfus2+fOR0pWwrINZ8034CSYKla8YZzGITSBJe5wWX6ObmSUZ+80ibdj0S9vLF9Ht
9bmmGqe8ziF1MhIIYh2yhRf+2KEygv6KSDJ+2XZMLvYEeU7XNZnz6e621KizK6n4AV+VsfEE+grS
dtGQ+hL2Vuy1dVSzdlZn2L6l+DSm1c6o8VEVxD3xtoD183igs11dq+asuxwkffpz3Em0CagOBTs2
kiPlWPAkgzI8YXVHHgW64bNe7JDU002DONJARpJ6R7fonW14k653vDeR1bSv+ZcIxLvIAciZCCCi
d5hHpRH6BnKrReVanYXrlZYjnSUX08gi4Tw1zJy5GSzlG3hZJnN6lIOZ+d4IDglGXJgvnR8VJSgN
GeOT063jlxRv5DIbgb7T+Vcb9O13E3PMX0EWlIAWCRklM671gkGDJCsAX6rirds9hiRQuuKI/9aT
Z567nu3h/08Z+gqZ0H15+KZR0wx554emS7G/7LUWaOyJ0k6wGTbkKhZttPzEm1a/xVu0YEM2TaNH
8hVdq+PMe2q7VcGF6KyLeVVywlVNQlsKOqjJcpcb3r+KskcMFteaNR/uz7Z+6b/dUCtwiHNjeiS3
lZU32VvmHVPuaku9274+x+vr3oFO9vnumtGrXJCWo/kjWhEmVIGmU+1s5DP3hHmhzSmE3lQpY9WE
ei4LXFd8ZLjPnDciYbdARjl6WapKun15gekcS9/bs3rJyHPvrwrGnoBXv7iz/MgaOm10T8TV6BQH
2HsAzWXvc6qmx0PbyHDRYJDtNPJ19dcnqmdp1DWrCLKK7uvFUNlmuwnQRqHSQx/Bc9x9lThS33ek
r+zUQNrj29B4VtRL+RFJUKoDxkigva/ymfKClgqg3GjWj+3WOytvEVIEpO7iSGvOXna6gWwBSEU+
ZG3bbcwkXPFp90kYBHNJ7S20fPicnH93n5Ok4W0WMYpC36UaEpyXECO8+snEaOzAQtWsLirQvm5n
UtSOV76QuDp9yI50QFQAXWlM/WjOamYTH4JxScAO71ajlj9QYexUkIPklaXG3r+4D0IRMXKylpA9
FDouwNb+6xcSZmgKddCLLhgDCggKYm00zF2W2oDQT78+aYHHi83yTU/D1QotAwV29sUg+K9OcX8o
hcexujM+ZyOviaTi/oQ+bgrYzqBtVc+O0lAb9eN7wzcu61/RJngjqg6HuZyXOZ5tG2stT8JZdKoK
7OsT+AGbIKMcC0Wy+Z44nvIibkqJ/04DkLB99xUozeOfKzAJpqKq8HptsAFy6F1Rjsx0cAfWf3Fd
E4WFhswHudKEeF3ZRUc8NIZ7Z4Vu4qwh+g4TJW65UxhaL28nv5uU2PTKFkWIsfGLW0cKrjBZcibw
gpADu3fTAZfU0opu+tAVEKuPkzyLqlZZ4rD36foKM+HUDXtjvOB1t+UImBLDDCnqO5bTT5P6c/Vx
cfVi794o2kBlxTMX54NKMlCnJcHXDnQ38JnajqKYryiSieWsbSNE9HddIbrvMDFMBRnJq4AU7wN/
rVUCJ9Y3axWl7bw9/P/IyuqJvXOKS6gVB9aNU9eT8TdJzKepac/Ple1reyLFGDmNzQZZ4SvRg8Q+
ghnLXwkbP0R5RLRRX27GBR1OOLzSybziZNeCQFl20TPlXW/aGNZZZJMluC32U26aYJLRdSxFmifj
y0JUhXqUEVG5CFFiAQjnWBscmXXlvoZXcLShSghA0YBThxc9yXiUKD50BNAaWcT/EKggMdcB3frD
wYXblKYnVB5UHp++oWIOcZQQaby1yD7/32bfOcHVirq+beh9Cb7Tr6eiWqX0lsCk+Vb8eZq+Q1z3
sUdKRykJI+Of7CtM8LmtBERI8I/rIozpRSRPJDCr3PydT963W9j6wodq5lGyX4SeOpu3ljES4PPV
plpXwusreoMIeeSmDB91SR1toOkM/TuSJ/UgWLb/BDT5p5LTyUgDpSSuLQjp8x2SrGdE4Bcpk+nG
usjcAH0VVWtDIdTQRS7ZI/TUxvPJReBWTDb/taI8BrpB1RpibyGn4PECmJtqiTghIKx0pQ/NiB1/
oFFxtlK3ocnIYitHbgjuXmb5CGBTQVY6FcdLh91meS5EqjHVk0ls0/c/pa9i9xPaHlVl/4W2Qi5Y
kfLsieGk79u1e1In/qaLCAMmPi/up2xwCNvwOkLrC9jLl6kOOND1vkpJ1AIVtdUbS1FTqNVrhCCR
DFyjq4ZUSDTSQ6ysRGGGjXTHLlP6I7lStwKFOvejrvd8FErUdbnt7NcgInv8uYReq7lxmZQy/xnQ
jLMwlSpdaiKziFo4KWnSQVJhqToj5dXDGKV+ZMRd2Sb8rntDWE2Sb/Q7f95EFXWupbynZx/wiuXF
EbFQBBFz+xX9posoZGGxFFzCjt5sM1ZedIAtp/WVwEFWfStedo5VunQUgMIJUbF6YWSjI4v9qafY
YTetTxZtlLdAJfGi1+9P6towVMKzXPH6JpttL+WHTMRGfptXPsQNVg7A81E2Feb5YExaqRPJcds0
WkXOQU6CSS8p96ZF2syHJHhLd1tt9W2H98ceZDRvZV0j0Irj4ymqlRNjBZwt7Hvp6xOlXN0nxW63
fUPxm4rU+VleN/p9cfLdpaD5W6xdc7tYQrSHvLLmFFaxVDVZpj8c+ZC6TTLa6qYWBx5jvYIar9BV
VbY9tbAVkXqTgrLH6weXty/P0hOnf4xkED/CP40OZ0vVqpmkOseSeJdiQkLTRbYxYTzdKidUgQ1j
Ii8ICdPQPtcmFszDKoJdxT6orhBjO9AwrdQRAqcGG96cJbf/muHZXQFbAPo7EPi7SlcNOEq7l8jr
cQBFmdgM+2BTDWc27jJsZg2TyCalFf+vjOJeMSkPKQjX3Nml2LgBjMap3F7+vUrIGpSuzD5IiXMW
/9ht9OfuNbwg0GRcuDCOSPtYwB0DswUFMgAuVByi9znWx8gWFYAqJrFTVrVfzRrCl4ZFnTaKuu2M
s/iOy/ypFwwrs1ocVGMPpwEciN45uRgo616Ngx2BauFLpwmo1PfiZJ+jNDrAS9jW6EHyJIiHxJLC
ICeOhRsUfCCmr18dsjvfhlIqgABoJrBSRxnZqP0iOWY6ZBb4MWs8Q7nZRp9pI5HYfT1PX7yMW7Rn
2w1PNGP0F4+wL1NJS+i2M04DfSsTkDoiSHvGXW3wrbTmv2QFksZIPRCEbcJLFlVeRDFKf4Gz54Xz
rjA1ds6X/po7tSfxw3/H/WTIdMTmaNH6BjoKKWtd+yQFo9txtHIi7crjtslnQfcG0Iw+eV369hHC
oakfg4hW8dVgZPKOtG6ilTdkzDSG90qk0Q4IlfOtiX9hhzKcqUK/+a2PrxXjTpi1vDAvvLzIY1F1
1+CxHnIAJDL8qhEysn1fVZIDcuBRtdqOgBYN+uaOG/Y8Kegs4hO9UaM4Xgt9QAKu8VUCQltA4oEU
iU9mvfyLukInjc0ef0wKB7Scvi0d3dZTbaOIFq2hTtbUT+aZbkBKK0DTn5K32YUwSOWoNcOtXHZV
sXZMIECuLj7fxsYRNnBLAWNqyCBP6/6c6gZMZ+Eyq4bFHSVZaCWYI9SLMRzXvy0GvpmHeSqols1w
wDZYZO6Ol0x15K1y87oZUcV92Zbn/iD7Uztx65cbURKTMtpFkTtc6ckkM5DyYOBTQlfg3SpRobCW
uI2BppsPnS07ZgyCQnSlTVolcQUApAPr+OBsYOl5bMG2ykCCBmnzpRspvjwaNDfYZiUkm9IGCjvv
F3aQsChgxRzqxpYnnMt0qaWxmLNaCNsinIykgBRSWfZgQgpiTbZOgI6XglEENcrC2aMxtPi8Jzvw
ps+PWFKSWsk6NvRjI10WZWny/exdZD8F3rvQ7gsDxKncaxj7IthLegR+bIgVpgNRiwhq1yj4zze/
tyvzmxn1pwydq8rRIPw4MWHI+s8JV1QRCxdxuGbvO2TC+kfjmumcjc0T3wVM4afkKQJT+91dB2No
XgEutNqXS453kjYF3rIpLRhob6JpufzHxVoj/6RwdxwgszwhlrJvZxd/Lc3+HslVPMnwxvqzkSME
OZyU8DssvcTT4BFkIjX909HOEX3cGsNnPAKBmwlu894xX4pg4lvb01wESDMqFNg+PRiOTRgOyBwk
UK5hv5ThobjkO2Xjlp8oM0v/pEgRr98BwZ+owuW8xlD8rSyzWIPVchxXVKR6P2t7w32lEwWFVSrw
Kybo5+OKAo8jevaSEMBhH6BCe7A9PYhbbymuYcFkjsABU2/XSSOJbQXQ950z8w2tucNXBIziWCFZ
0hNc3m5YoIPGnx0oOlgeLtJulikZXuqh4vRYXzUS5Q+Ha5yP+SNM1cL/ZU00DoPYCQXQL47LAFku
B8hUyRrxAc3IfJWDXFWCgkoDU/Th5cgDtJQaobiRKTfAvkgviET0ZfY9NtpXDhck0xgnuBMtfgn2
pOqSFx1if8Gm7e5rDt0An8/pbbVj9lqoFLDgGyiOCrJqI29I2wQER/KETHzIrD7e/NQL9eP5xxfY
yvuFQc/FvxGuH3o6qI4KDwfGreyz3yOrP6FUzT4S0nwPZxGtWDGLk53oVrTIk/5ExQJgeLXHy7lA
bJmo3ZWmw9dEz3cHWy5opm6YMKUh6dvjCC/JfowwYoHr5HZDTYpqSkrhMYBumRPt0M7Ea27XxPzO
v6yrOXsoXVOIXU9wIeZE+25bw6atYDcI4LP7xsbDFVdxaq91Jsli56K45Hvhk9EOpKPANUa/XG1u
Ev+5Y3PPV79cZH3Ne2kNE6/gJ2QeCODTMWcMPEJtir699FL2XBpT2qQExQS8NNidYzIumpHTmnNT
kLp0hjP3wvGRgSoKpMkdEpe2/yH8qjmM0WJZ5ITrWwHAdFxGdTUB2InE+bmfcV8xSG2xhdpvMOx8
5onUzzF0763/8VU1e/1uBFV+znc/2tjeL0OszyyrUCmJM8+JLjFi7uBO81dY5AmVwt/C7YqwXVAr
v7wHfkJDnTM2O0XQDv9o0FbipiYmKBqcnDf5UmjuWV2WxUdFutIodCdkiKjw0puDeEMdMLXsR1Nt
QQuV4xVJp1keHqWFnz2whVyYoROKIv+brJYZdQGlGglGAVhed0a9FNxaWvrNnwK3JEQKFoPMY8gP
11mJEr4TErS+I/xg4h5OjHONowVEL8YrtLV+rJFNxkmXN1ca7uJNXNoxT9YEHSDjaqk5NZGmfmpl
yI5VqaW7ZWO8BTVYEdsdwmAV8JeK1M6UfjklxORdNoc3qxlhYsEoiDcp3tPSvo8IZQ4+nXgpCxy8
2xvrNI5/rWnMNINcaLDDl9v7rSKqrBlFO4u5r+Uw/iXUvFIQlEn/qyPEN5nnvdUr7eLZpNK0Y7sj
WIjk3+QpcxF5YoM8q+JSC+KOpxC8My/bgmHEem3peeHAqP0p1de0rMbpfX68rUIuijj4W1VZpFEn
b0ngs7b67JF04FR1E9rqdIeJw7Mj8n/7gTUz5sXdDV6/syUy4loLdEpMVGpPAiohi0MSejNjIxrw
wL3mn0j3odetGeCUl/Sp/VfIisavRY2tWCCbUE4UhULKV9kDCsTOQdYrmK45dPUp2+dVGucoa1X7
kVCHss8DkjUwJKpR8Ij1nbRhjB4rDK83oO/l42kXnSkt5veP74ZEMKE8D3J3Dpz4t215ZPeS3ifj
Rux2j1WjsSzqA/aqIKpyf+kF+RKKrOe1TdCoZ5mDe3QPAsiscgWT+C+cyCKduk/DphHH2ErpK8DD
ahuBB1Waul1RsWHw0MZtOjheTGXvpEkYts75Iv9fK+4pnh3pVzHM4IV3dl05V/LVySpt821cheAJ
9MsNbG4PuAWBwazXOpCFKg1vxjS0+i19EZCeqYmsv4XK34hDKW2wD0+6TIxzXleqGrkCVvBc2ZNW
HAjwNS8YFxZE1oA0jESwi/Xmq7vbpeLKzMI5wADgFgX0ukn6a73I+TTYYA6QFRmU9uD1QBotDQe0
qKbgAIaz6oglCG0oHw8aDRn2BxcDTwO+8XG/yCUIin2N0mENc5LgxJG64Joxeb4Hvb5GV4Wrg20d
xYaQ2Bu/Q5Z96sxxAZ4h/P5TGzq7IzLDV5qWU3nTtovmg2Ike7Wovf/PGmr6J5Xjh5gTu1PtEZ36
Rik7MwWnrloOKWXKey8EWOdIzY1WyU5xVJp/T3Don4AU9XB9GjF4B9dctKXjDfiZa+cQkYPS3Fg/
XThLuO/k1N/Vihp0mj6M4lwFnSQmfXoo6rRC2bR25mV7SHXbWpOrxyovuQwqZV/plNE6Y2g4d9rR
mDkGbp9IsZcaSmjk9zgZIrbvTm/wfvcKhbK6upxFUYpxvoTwV7YvQQZmdkMg5LAYWg0hlc5V742F
6oXp+6Km2+Pot9bIQ1572AgsJzWi2A7cd6UFV3k8VgCLlvlXh69u+2rn0rz3PuMv5CAsOHaCNGRo
ZUGygFU7iEswQJ7QoMHYJ66ocgUCNhjq0++pNhXoJNxrTf8XYXY+VYuhO3UPlajjBp14uDeSH9YY
bX5qdrIHCKlaD3pnvflRRxRrldvYw97EBB1rfeY1uHa2W8xPUzEeIhJWSOzeVIXyNBCZblSijwN5
cnyxXj6dvWwiITMb6ByHu4xftirS/IP/4p/Tlmy7o/m5Uhzs5XHUJ6rPiZcXsLx/9VeIck2Zrepc
+PbVo41fXeJw6JCt+QIEDZONJ2/jLVL8s3IYkSvfp0GhNj4lRFj/iHL87RSNqwNgBksce0Nmay1r
rsg9f+TnX3OTqqZ2lz44OYuVMcq6+XfUAsDKqs/uHng2CKONmMj7y4LtfcfcgsNvvWhvy8vgDnWb
JuS+gbwbecUilsE4nSZq6spMKFaZW1CYmEudTCTwPKyDhugyUUFjpdxkrpSTuwvVyiyMCPkEfkD6
GTvYS+vfKWgVGtq9mZdMSB23LU43hraWv1tBZSzuKRWLo0Ky3DY+MUZ5Vy5Tds56HOIuYx5F19m3
Voh+S5Xg1WQmp99ykebQphomBSD+BCYXwJXyW4Rh54v22ywmETY0mtF4k2q+v7gXCRvddlP0Ztt+
duYAOlR+ijcA61YTDetcP5t+COnloLtq4PjXEJaiJ3LYnJ3Ji+dP1kcLuVekAXBB8xmVm8ZsZphS
H/o3joVdxkO04K9QNOBBw6ayvQtduGF6/aaQ7yONYyNTPhyjvxWCRi7QlI0EdQySiFrNvUSUuiia
B3hVyiiVwo49vNW0WBpbM/q016NkXS/a/u22V5RcfjK5/k5nU1oRg+XVhULcYZ6GkmJNlCQDPxxZ
/Z5cWZR5f7DtMQzr+3RcMytud9Jsv9w1DGwt7X+P3zQb5LT1OSy7AVbXk51pGS8GxD2zxTqmp4QM
ZxBrDfcCCSyscOKHTVLHuwWuycX22mnAyp6LQjkWj7ClwzYQ4hMLhTVIzxy8vyMNHrkknGG/1lMx
hWb3ceWc8Usy5o8XQbB3RenhVUUIC3XpRJgLGIaiwU+FZHCSuey4NnqGJ6qnKx+ew+dcZqlXIPs/
Rn/IpNgxunUsJDTDQ2OFdaIbjFagCBBIRcXn0QtQslxhmmoxCELtiwmea0d4TUHwhG46kUiVsxo8
q8sn6GJtRzcPEzmtFOavrQUjqQsW94xSEhqzf76CafDwllvJu1cRIThNYXw64uU0mP3lOKtqpdoP
Cif5+mGojnbKY1jAsKe/SqWhZyUk9+16Pi3kX7rCkQI7/umkx2DRV1XCPLLdQGMWNcsHYKvUTctp
1IINYfvQxWmwE8ez/ZZyxU4Lp8GFgPJEzhpxlnPHrOoDZZUTHzcxvJYcv78ULW/iREhAloI+LcNg
NrK4tJHPDYpRsTJrTgIuneIrlOYHrvJlwuSqzLE2UziaN/eCMR3Y/kW7ZKZgqRQfxoo3RGbBaM9C
UEU43bKNF2zsHALZ8gTv6E6USgkGN3D6RkFeOflKm52pNdiS2U1UP0RlcSVoKuGItESbl89XWyQu
rYEX5V+s1OD3iX5Z9aF9C6/7jgJ2iguMi9bhHxwea5Shh9tB0Cw9odNy4Wt7xkVeI5cQ7CEH99Wb
6aYv00/pB/hm4mnUaFB/jW+RAvM8l9BHh5toFF3HxBBg5n5Llx5xW+aF2hNjcxvId/TKHla5ehh9
yg8ua1odAJHCRlA0HG0tCoBBf3VXx+ys5insqthJtF1XyWqqJY/7VkhO0So75vExdJrxTwQFGYQy
S66pI0i6UowbxFCZ4hfVSmSYqzcmevRjdynygu/3wVRnKydZL123XUxWOd9RGyKzabmbBz+mZPed
cJo35JFlniBHZQsE/zmLlD0msA08/HWFjSq35FYKWQhnH03dJg9vbIEnXHjHywQ3MPTCdpdWgX2+
S3C4hp1d+14jhN2E9YGadDS7Ht2ppG2BYwLz4pzFKL8cNyYUBipF0sesGzEcCo21wt1oarLTMFEa
dy+xhAVY9egl4TMWHlIE0iSZ8LZ2YkWFmZkTdRfS+f4q8P1BpKdiSB+n0b/lY5luXfRO20flUaUZ
bcJEgpEzSRl69mnH4HaPLKejgpLjGWU1pf+Ge8CMbKRKAq/+k65Aelp6i2NuDPQZ7MPK/Uo1PbJ3
wjwObJbsOcw0W6FQiJhz0G0WPwiUq0ssjtPc1Afi07mRiFOpUCe/djKjPdzRUyfVklJOtLL2xRIE
a95NORPfzzlqkJlgVOdLP/mrcEiLpYBkXNioIGaJq8CsNg8DS/xKDp7WaoFIqo9bH5mrKhH8mC1K
p1FRsuEbLx0h8sAf3+MMN968rDnx7LcfFCcXEBxAZoyRvy7enI0a55Cnax9ZsrA9U2XVDi8mR5L5
p13O9qopR46coq3qffovFMB7yZijvbpUK3Jh8l5IcX1mj9R0DDLkL3U0ebm0a3FzBbaun/WNEk4A
dmsg0BcAXduJrYSjTQNuoQbNlCSa8RkxHVchWrRC/K19CIfVt+TRC9sKUIJItal5Fai4n4u+1/rw
7IWrDw8YshdW2za9TjfYSPgL6yT8ijeU7YQHld41EC6E3GR6hFvOqJ1BW7m81wty7YvAF58bAv5T
J9Tw7thC3yoh6dpC1jRm/hD200AVYHKZi1Bs592WOYB9yJIxp8AE8YuimF03hRAElT4k/NvAUSuS
vwMCkJmuZ6eTbLKw7M1zJ3OP94Jlj0lowYBvaTIp5zxsVb+es+/w4VnrU0RpTub2OA3y7YoN9R4r
gS0nOtHdIoMbSWZ5sCNuoYtt2Eb5LyQyPEQCEAQs5TTbCAW9I8N164ldCx0IEldYej8CHeEdwUBW
WGKGqghk06aCUH0ZmwfKDoFSJMesdrA+1fEW2l6AXEDGTOF6QDru9W01gX43NiaATKo6PRaC36ld
4ta8tuHUd4XnH9mZuTWigfB1AuYQDbn2nqFZz329ZNwSZ/ivZ/Gm8WUbnKg5Dy7ySQDoGsGmYi+M
65B0Eeo1Agxb/QhD6w2EQ3GbOZg7/UGsAU7REf8Pmt2/Avhz9tQBuSZSMoLH8ogcu4DmSipanLlz
Wwb+NEN5Z05b97cxlHOGzI6uniqoyWvKeK/Qw5MKIa/3jlEts9vGS3cWIlwwFr3/Fo0HZ5ePsJUR
RLCLzVD1aRqbpevxfg8s0Qc08FvSF3OBkiqOl3ox8gW9PdpI32UCNEBsfcwPY3DV4cAZHEhFi6nm
TJL7dXtUyv2/xsRnsLAIwqjhEl55ZrEFrvQE/xVSabcaOjhPPZFwKn7gji1WQXUc8h+gxyngXrAY
WjOUwjDPqglID1meh7ilbRKUuK9SWjQrnCqQoS/JUWglvVZ548PqUXe+pYCwVSQHA1oIOG236p/a
zpJa7VJctkXIDSwX74NBlMEOkJ9aSLGfT5oQ2DYkLy5xb51MwUzAK5K+ZazcSCJhAX32Funnqdpy
5IEQwmAPmN7CGRtZMDzFOHiY0KcN+iqrDa1aH12Q2ZccXHUruc9apWJ29lCFq5KFBPrwbJSMqbvT
jpSSlotVWj5zkQMlT/tcnim1/xOu5Th4kIUaELR7icEs7MpRQ5c8KvX2+cDcWG5ZL0Yr2HVqWl+W
m4wezYjOtgDbG4uPPnsEVsQj/2vEHLTqzcNmjaTIk5xqI4+e7rfUKfti/0pLXawqMkFPLABLEtWE
EmtSpC0vPmnsxE9OaQE/5qKzrJh48zH7CleTaisen+osRCHpu4x9ORVDRIEqgRX3F3DJgsSaV24A
7HlHAPSzBGCXqBYJqlD62wdA3AFZC84kW2blxSgx6ItaOrCt3i4l2veufsux4ZK+g8BR9sN9IigZ
TEIzdoGUMq5fp7fWzXPFybizMLhK4WNMb9Mgway4LPWMOFiu70N9RKyMGQHBz7FFGlsWD/JzvW3H
HNxUS0iJinydM4LFnfQZUrnVOLukxgn4kB3c7xRdUoKTw1HAQTfsmwLpOyyvbRETKTXPY7GbqxWT
8kw1eXWFBCpbyvZxcFhZoLWEQgfdpsuRQlUS/29A4YqqMSGvPf82nLVSxGcqEPWT9Y6WkI5HkK4m
nq0JnHkjR2bnXKtS0QM0V36JmRqYpTEjSqwG9OsCZDG8YgUA4x37mX3ZtZd9fJwluI6r/uuDpRFv
O3/eRlzG0eurEbgWDiTJzrquc9noO4l8lXHx632IXufTql6elNdDkVjrBb052bdxo9Qx7tEuwIjP
ymnJFlTimaLUBgSbZ9PGlOvbl05+F6BctIwGNTuoLMrMVNwKjcOQOmu+YzSutdG/Ldmpi5H9Yha2
4p7/UFYKdowf9gOHFT+BzpSGxLTTAHoSSrCOk4mxtHqUU+PtLDdfK/sh6ar3KzbNpRHmD1RPt+YA
Iz28aicgPFQX04WU0W7ux1TWmsuSUA1d8k6nIrXaFHZTb9yk8qAlLm8SckAZSi3ZNyCOZMFwEic8
mJ8lS5Clsr6+1N9rfHN+uTSd311WZra+N4gHTewnPs0AFMCBiTGx3mXWvU1l7YmgANovSDIFJSjd
oyL+F2/T/0EG42iN4r88lM4ycL8vvmfaqs64JFqJRr0iRX8hhmgvBtt+zS7np3ZY5jHtlSK4Fvig
cEetWJSxYQVDz62W5hdrBG4yI4YZoZtrGLUZgyoKs3csHm+sRl+Hx5ES6ddp87tEB1iTMluWVGHc
TktPWgl2ZlzBc8rBGN1HpF6keNmrCVQgm7zqZgFd6JftaEZn8OAcdnl7JKy/08vVGzgh4VdbYrd1
snsmkmXO3/vN8zThpVUizGORz8xncxkOAvghhxDEWwC3EgoJeZA4SxTeX9VmXIDjvfXlWcs8Fqxo
5v7eVm0MiXKAAN+B6cwHoTjQhqWoGt3tZS7Rv7nDwz+alW6NVHmy7Boc/PO/PqYjpwAtszyJo/ju
E5+8sZk3EAiOtoaHv5+oMGVa8cG8hviIgla3lQUbfsuQul/la25bITGixjjXexxKgZLoHddvc09m
GK4iD/jCx3rOgILGdBDc1MQy4TljEP3PauRuhLTP/HGTK1vzZ6R/x1/aBncoy2pz7NHSRRmLywh7
o8aMcxd8v8tBX55+m86ekQsRCPAZpsanmcb/oMxMEijPfq7zaToEzo7Z2ucMv8d1Xy7XM8nQYqsF
5GC7CrjkZu0U4qHS+2OQCuShv3yPnMCcrlRSL5y761Of/FyrH845Wbhbt6gUt8IRahaI01ZR8PFb
yGmY9iQroPX6bkqHxiiBQHGnw7ahtweUP52/InCUADGSpi7buxd9i7g4VWrTMYg6Fbc7E5vLOSEq
AynHszK8HskksPFkBzaeOW7WaYe3+OJ1u4dzrWOEX/ang2SJNPgFAexsiIvuK4oyPvrlruWb1nPk
DwmnrgNLWcJTNHbrXoo9sdka2IJvJ5sj4SJxwxBxnYaZox544OYNI41lKi5pEto6Y3I+DO5l3yO4
RiC076SS3DGfKUdPex+/XoNcpeTowdID6M8H3CQdU3brVMa1QX5ngw9qamyMkYVy2FxpMupzgUmh
Cieqc7CkwXa0h8dHtjQ/dFxvFJTf/Hffm5HL51vD825Hr0pkc2iQ59fQWGpl5GOeYGJ4RXI7IWyT
/ms8d/o+D9lg0/+gM90U5LskCCkmuwtF1mCRmXzRjZ/Ip4Mj9Y/rF6xOd8EOsTZX+QEge+IvS/ni
Hu3pfVs2G8ppZiYJBhexp/JWC71oPBZHD1zAdsPCYjVbmnSLJwmpu/ePzgUzXTnbl7ja2co9A1ER
oUhImTM1lwBJypG9Whfy1WSAG2acPBrM4bMR3hxOhjm4R5ZOIFQZuFBWm7y0xO1q/BhIWJaf717M
5At32zNMmiwe8f9izz8aj52gLBZ4NaMEoVsfQj3R4OwXa3+jQ7Sf+S9LFuYFRl7txQ5GRs/jHVAB
AzXrCw0IFV/UA6cLWdKEYHIQ77QlQp6lGernYukvOaWco3OEqcnJlvEbm4x+HpIKh/S459Ui/jK1
PThlPpBuM+dxKNTecTCdez3aZ1yfGiA3NYEg2oiTqzD7YbZzXiJWd8HMkSA/f+KIlOTVN3AWhahl
L1U0G3VAYBhp9Ua1g3KT/wChPhHaPH67aaNBaGxlRFkt4skMnKiThno+crQPz7F4rYIzC/vjqNMB
RAf09L3qjw7IpBUGVCHw8bbd7tPPoqpF10OW0/DCz5HrErwv0in7yO/xmPFZ0TstpfyuYIEb61M+
PBISx8uUJFtMbOSMH4FcCvpeny4AaABbi4tcHyIwH4F/3dN3oXIyRNsFjYBcdbLXvCgFfkms3lS7
Pb6mH6UYzcUpBujbrfC0GEnmOhARchYejKujXALSs7dkggBa+3mpPfiJbLQU83DGbSjaBmSeijW3
8S16weBIcyWlGGnuOAeUY0mK4qe/M+DzXzDxMcXiAhN/I9o92x38VuVd+GwRjbuOxfW8Jgo5ZfUY
lheaDBOthkbTyHurnP5QRNsKzeJpyjujGC90q0T2Vfx0OnT90iCfApv1GBYF2YQ5+fIKIolnCw8o
OgwvkQGKl7kxrsY+SucVkHoOdCT3oMqLh3GRGK4kqR1/vlWLbqtEhsQ4MAo9ryAJoFpp7XGHq6Xp
p5yC+EQAaQjrQV7AMTcrYL/3izRbeTkMAFpsn5k9EtIlkjiXGY5D8OsfV6JbV0pfLr9492dWRBXu
V9Sf+cKfLhqCEiS70bUQ6/drFlJkddKp+9OpPICGdWWdkrhjX8MJcC4c3UMgZRFPCZxzYNycrlMX
woHSXbAd7d4TROEUhporgBBv4WIxo9UUirtW06GOiLkXXqd8UtZ5m2JEbEdIH5VQGRF2zWSJMjoK
D2pnUQaQUfwVpML+80nsEaOuPuaaUBr9t0VeZ1kBRi0aHj7r9GJwqV6dLz8mNNZ9klt2ANkF5nr5
zMhYAPBc/lBh8b5RrlqFZ3+mZmAZKFRgLV9TrjTYRyDJe6SDLvSUxXkTg9xF+/jlgaiQ/bPMn0lI
uOONtX0lO9Z3LZ6ArDAId6ONLtJtHcomy01lW74+fV7hGuz2b0wlcLTcrYOOjvk7t2KJGtI4VYPL
RQncfi2jhk+OcXZw0YTc/+jSfsaIbveMyofSRJ2rw2/SpRv6+h35JIvwl4IoE9w4p0CgvHDW79jt
Ts2IsmR5pzZ+oJy6r6cTwJIkBCWVH5yTWaH643mv0e/vd4djnB7pIazlItVpohb8vTT9iZa7TzhC
IcnVxBa2BXCRZexFs0vNZcOtHPQ3PE6zxnPt4OjRl9tXfS8TAkfkfQRp4Fir3k/GIOwyCRBdLBly
HSs/M7S7W2hKzCQ3gd7k3aIXiNc7YgZ1GKcbd5uaTnEumphRcNao/TKjfkgZTlrGS+xr9c/C2l6X
UsHU4WOj1YyGuLR6/TUaLcwmaRtfz6wVfAds2EIUyJGNStbLoaOB9kiUx+DBYZA4VLG+5miOD8Mt
1clB1Hk5xbt5+DEvWdgpr5sKhkjlIWFiGtiexlZqt+rxNAS47HrKxbS5Z0/QCq+P53vZY707vLHr
KmU49Yf5pA4hUHWXzhADYL0E55A5BmIA55hXb932jOLbiz5vPTj4erhQjxj1QWSKPKNKpZm+GmLy
4Bz2FQGV4FoMUumEimrySfg68xxT0Y205SBoNkfj7DvPyWdw0EN1KaHvQ/2aOGkAGxp1zhNxFiIq
BoJRlUrfez1aDi8hvahdtRyIosDpdjTtU8AxIvQ/Pw4uow9RL7+EnQEQg0zwJMV3sRffx50RBtdH
QIkepoRZUIYz3Aq32jQ739k1StO9z2032y4NTR0qCPGb+vlthuMXZ2MNPK4Ak8mw8nTpmTvaI/kO
dFweXA6Q+QaxDagS+x7Hd8uQHonwbFAYvrrk0QL2nFckZdbeLrSX3KGf9QPANWBLOo0XY/jlwQme
WhaeTy18JMhr6QO5ZrwVGrKrAb25jDvPS71Ve4hRGVcYs0lI0JWdp3BDrUtwILTNakdrrMNPVVRP
ODTdsPyqF2MjV8MftkAfVay8r4XQ1vJERylljTMR3OP2Zdtj6nnjy1ccn++m0c77iiHaLWo9kn5l
9RYvSCeselYOaZAXp51P2+NwkIPYjJN6a9HeKUIJwSnMtGWorATlQitSLM4/IKTH8Gz7mbAo3y2k
PkP1kbwnAcMIJcoXeiLEkkQCctb+mmLorwhzT/YVFctX5XVMox8E7Mib4kpk6th4h0LWeb0BB37l
41DVD6x4hLeArcFjs2VMhul9rAeeJZXA2+Ik4TE4QZnFubCuAxA1Q+5WxkR8xEOEDCZMz0Z6dI1q
0JEWeRpt5xJJFxW+BQ8Za31D6iuvzhqlMeZaqB+2/nrW8zmPrj49l1249vrwPiaOE4AmGLFP6US8
lU0Dr6AZ1kIBlihNw/SzyHs3ciOcM7f/mCe2FbBZGow73cST6gW5RpCgI+YLlavABgUgwzhD4SzT
XecsHbZ7fcEcU7uTXtEbPRus+pJne5JS8FKPPEnXxjWqWgWCgEMnaUo+ta9YtIS+tAKMk+8/ER0n
FNqOZakrQ9Ou47jaEE4HROIIxPDE8ahEYLk6iefe/kndtNLERPs71YTtU2fxx5MCjXxL/DwUMe2y
5SasexACxD5aNTZtqnE4bn6qqvfZMCVO59t+su8usAy8YqrNA6dfIXCqvpfPzVXXP1DRvnHt9eKn
YKkLId0SCo1vN8F/UjpxM16OH1/KYFKjFzcsv8BUu9qZq13SpzpMPDiOAkMNrOWpcvPrkRBYL/3B
OXB3uKBpSZUWPivLUagtlyC6zq+pSzb3a6toTeVLWoq7mhF99hRBAj7jizLrCFlqa/9HjmchywjE
GM16DeLWv/OT+Ri8O5YFic/qbED6+nkVcJY11790oVRByI8zYcGa9gtaYvEBcYgIENhHoW5Vut9p
SYmQ3g9SJI7hRnX2vF4BlwSMjLBEzBq3FmV8JmSqjyjM28Nb5HxkBkOp/Y2uypF7GqLFUOICRNoA
hAn71+k79OBEgn9mQDVFZ3sNkB9RSZHh6hI/f7oi/OPTmXHNcdfrEvLH2Fu5M0nEZPCaKBRqfh30
mMo+POMHQVelJ7BUFHNqrRUwNKugDPXAY91EWlDtJEd8SFbIyUDu6FecpQf5fgASBZCcTruHV/U1
W6Ibuk7BJ12OCvgh4KRkCw0XDoQncCs0w79Fwoongm8XAVHGPF0zjddXMcj4mVncdQR5Nw7SsYuA
8hyjNaIGsjN++iY9ibRwezOWQaSy0trJBMCfGt0c5QyVjhbQZW2EPIsBCtVqpUnxQeD4fo0dzt+X
7dxiHePd1Zv7MQ5vRijJ0YQLXnmTg6IA9zdqnkydKFDkz2AXk4qjac/7i3KBU9+wB8f28pVsv0qj
R8rBz2U0zrcV7c10H714Y0TeURgrfN4a6EdcptwNQZQAc3RFnQHu56usVXlkUFBPML8UcN6IOx/3
NzwD2otirSdx7nlpfbUzmkJXVTvZhFUXLukulA7mdfBIS23A9t+ryWQ9EHhYn68FK9zwxrpD4bIZ
JLYycwWMWfJU4hVvn68Eya8GPfbIVIFZs3o5MVaYS1Xnx+gmnAMk4sx84hse0l1ULsCg32Te8FGY
Mvc3kNe4eq48qL4UCvOFoNmrwggOoVYMedRxMqcfSGTc4IUannwTOCEuOGPjrapGjg1/ZnC8fQtX
3YL43mWK48aegJOyjMwCAsV4W33V0E+ojddZ+1XIDlhFs6i2ecx3LdlIx7P5YWMAwgtbMa6mu/KO
FEmLFewW66G+FH7Q5cXDnysbve3Z2Aa2IuuQyjLFTP4s/W0WDqPQkGxpg1A59IKHHmLQ1JwHWdRQ
prtsdCmft0Rjy8mRDbCnTKJQHftBOHWlpRZKwtJbvW5VnaOTa6AH0zDtox864J5rqfqJtXzdj1Ld
Bpnm5f8886+OF3LVnaMM4fEaX4dck6PU6ncTAepDFdf1l2BPHs+AD6FPjt3aWfY5LiAt7ham+zIn
cBfvdHHkMzQ6SAddIOq3+DdLDRhr0qWMF5IAOr7VheT+/xBJrZFmcMQtpiV2mkTcLsgV2eklDYe5
cSL3gqT4AHaRHjdd231h7T5jMWfQkoCmb62mmpVpPQnefWi8Ix/AINo+AxLIXwMXCkZNiHaQygQR
SxcOXq22CONQKdXev080syDuo48B/ATjVyDQKpzwOVdqmjKs0HOZ3e8CY/IGcf7ZByaHIpF1TmSO
8lBKVMjbBXnYkxVn6TH8hXLf85O5BKhveacbaOP3cgzCGQFlrOWmP5ucARPWJwFPNvoL4dKNRYkr
Z1rH6otX9ZNfKx5Zk8pxJTqxAiqR4gMMiuuNARWsmC8O17LzCR7tmoSo4rKxgEuNeeL+U0OOpQ2k
gAEO+Da/M+ww00NHVSwlTbHp2O6HPeamz4i/BdXAak8zcN+ISL+qX/fyy+olZNzVqHs0noVz59ND
wCTgG24j3wViXCYofijRVceU96Ub8Nm27BAyCRfCwDmknLtOCO9Kw8NBeml3uto8iP01ACRhBIPO
Xv37h26u0Z2yB9KIF0R4NI+b48f2esht2RniCxnZ7st1dMBAyE89BTs4odWahlBniEjLEKJ+xMkV
0+SaRQuoaly1WPMTHz32mdAFBuTAcXYaqtngA/ffHHHjontKjqlL3pwk52g8JBqdB9R0VmCpnafq
o7RKLIfjmbjssk4B7yGkcoK+5nS+PYn+K18CJ5UCAuMD5crqoaZkmjfkynKwWwIjMskHuJS5etmU
12kN0C/xX4c8iBRfATl+1N49f4EAfvejnrCQ9RYos7DQGFdA2jfUxM1zdsx4r3xYH25492p1jQEw
zyr9lHRGUdMz89dYGUHT0JwGPtRmz9hoUfCyLYt80C0GLxf0aZB94IXzT39JGQ1UsbCSEaHiZh97
b9b5FDixAmBUwwNubDXBcXK+8+6Jo9cjwmnlFr8ygOwwUXC4sOFOPp7H1ADsfmdPZkpsJQO8RwWK
Qjvwt8ZTOU7g+TP2OW7042U6l4RRfpG7tBi3fh9mmCVfJhmw6+mptcdUZGeab59LoeJYlZk1xFWJ
5C7xOFWXeT3c7c76jCxk3NwZFijE24oGWd6LvzbIOI7lAelAGeQvVIsC0eLUBaue3USoTbCIDhU2
tV+g+BtLY9imzYM5frs0yROQlse5VySVHol3rL/wYtUiyxFY7VkTMYaw6gLs/Q1gutqD9JqhlEy2
5DCJyc7fFQxRm1r0KP3+s3ZY+SFi6FuMkaX9vvaVu5zsXgiI+kxxxkAg1JLWa+OZf3LuOtCu5TqG
yMJH/e7Okt0y4A7C3JHVc/fM/bBKtZU3M26kTkipHQIILX+5AH+uS0LeOOZB0F8aOC+ZrkYzQzXA
BMhkrsuYVczzoHu6eINwD3i/Yh0ASjno9qpea8JU4sx3zlCfRyI1CcqyXwXBrkIqSx8BIJ0PvjgC
Ob0Cn78ugYGOTPInSk+CuqBJzyXOQy7jM8dU9Xv9xfLzX2Vy7bh1S4USrcrKwRFksgNio7RSnBOG
jDVJ7Gq7fgNTYHlXhNVVk/BFhXtCcndZpy22hba6JWizy1GCQ/mKXKuScBSWoTXX9lXajcw0ZwvL
T7sJMgivyg+gvBMyLweg9Lkm6F6XjbhNJwMtDHAp9UsfXm0zl6LFon54qqjxZbYLPp7afS+wYXRf
UjCzBIacWdK0KZItTbLlv4FdqnWR/iQ1tsP5bfw4T2msHNY0VCn+HSt34FAndfj51188uwWiJlgf
zseJgREcelp3K6gfurvAgvE4GfM3wvk+RRDhbvm+dZQy2jDvq/cnS7ZuQEH93cA8O+jEHZirNHji
R4ffISVBkoIYD4d8n83T/eHUXlqKx5v+Vha7/NuYAEnQONeTAifr3mRqSvre93S6jQOkV5sLjxfH
Zy1nywDC9SUeZn16/TWZ8DmIaGNq6lSirKs9k6xszmp0GZXXJRYNslRd15D4vFfqonqyWZbhfnEF
BNFhf8ntCjbKJEvw5nM0ZlR9y9HIWDytcX7DwQVIJgBo3b4pgvhZz45LL45P3i0Uelj1N4AmTfxO
XXpDiAjABMsyYzoEFDl6UbRnXrubaFIhEHiRUGwp5s1A5hhT9aX3W+qZ7igOWc2BFz1XQcXazVFG
pXYU66nM3xwdDsdqhlKLircTjxAVhiBFDavC+HKLpzZqp50GjaCI7UkJJemKE33CX6m3IiWrbNug
9ROons5JcNamvCMdC7wPPU3X5bqTIbrsn8QNsThfGy1bHkq1hcB1M3OtTQfLIBZmHp7GmRsN5P56
PCOXk6uXxdUiuLdBcO4GOi//xsa1wUk/tGy3jqNF6fcFASfvGQHeN16IA6jdXjFohW61LuBWHbxv
4aZopVWm9jT+ngyo7lI2WFuJVDlYvknLyyZ523NWFGneo5KYvhipGp6xdGy2a4z326zCU3kt3qF2
6/Zi+jAw6t8tKtOMnVHF7kMGfvTOkUD5uXydw0MYIciHFUdi8Onlmxhz3rqtB93WablSWBsVy2JN
n2rMWDDbiQcfHzlI68XAv5uaTl9mGXtde7a7TLKF23OJHz+Pu7r56nzpH/Moo4rYUzLQhb9IkEWP
6FvR73altSw9mGur95RhNKEH/VhKo5TMsH872vfwqxCqQIkcSrac0BBFFXm/rCSG1ug3lX8+zJoj
JKH4UcUSjd4sZ33n3xCrphdcONPnlbj8e7S3OzGDQvY0VKqkb/GDHQuM/TYSwCq9pvfWIPUjEucb
n4nENgeC6M8Cwqz1FOX6xe+S5QU8HyT+95HpG8VzeUlbF0JcKB+ncA1WssysaRkotQtFFE2z2k6n
SRnVRpGgi8sG4aGcuPRPFgNOz+e2A4UZQxrRWWXoS+TKEPS7z6WRxTt9O5AQYhPo+7v+Z4XX5qVU
/XibCB8DHlQAazIYlp7HSbDjIc6CtvK6JBQcleHNu2JJ/5kxH2RBi1ElitrMMwDuo+hZv9rpH5m6
5rF/QpW9o69isVAEmvRcCdKh6NE90obimhx7xuhc187knbWjQXvG8UZrRVWFUWhZRV27GGA9Kx6f
ZUD5w8/Cr/5XrIEqWaTDGuNeDZnkEEYwxYtB085y4JU9BG9/ejnkmleIwlZB/FqY/uN52FRPlciZ
18DjyhszDGc+4YWYZqexGeEkRH82K8NnqxtsKOCj0oFccC4ALHM5pSH1GsXZhzg6CYCIsK2/oFNR
dHlKEv7BUwbQ0cf9PMLgtjZ/WcDwC29PTPMSTiFpd7FcW0gaeUSUV0rQGbLfSuVTqldDZ3m48est
rymPHrtTROZoGmjfaosDjgqj1N5o/+XOMNnvgOy4C4dDjZpd9K7jneqCRPXt2UmROfWI655/s1e0
N+W422EvKUVMIUDt7ZER4DoiYgFJ0x/XUCEQJeBwaVx0Ax1jUX615d1/z9iP5NdcW+DALfmUBwM4
hlSGvU6sQ/h8GhmyJa2Ja2EfkhO43KfT9JcRjvPrOP+6qoE4S0SJQCGGm1Ig3zhfVs6F1LYmJoEH
gjPvabZTLTcKYG8TzbUrVJee4H8v/q5cJLLrDM4CqnAhjacsiyRhAKX25dcUD0VlCIzjfkfgwVbW
2rDDT1dY+1TP08XfCRGoaKXP6wrLn9k3Ge6/hpxy305orheqAvXGqIBqzglqtUGCPWy1T+EOO5uA
ZG7EcJUHujkS7kMp/oSYhc5faIu7oIS7VROfCZDXxEPTelyLuuLdcqRqC1IaU0DMtdJhfThmQMZf
ezYFLjDWd2VHwL6nDa5xx/JgyVRgKr42rrV67GLSidmukavWx+6SO65t7vnO5BN2NoRNOWjzrRdl
jHpCvYI0sbDm0bsBgf7dZaI2Yfdhb2GStSKKmn7e3JJdeaGQL6woklRxwL5EZ9TvVxkDWyHs42rZ
n+mVYVF4grGbrurCpGeZ6AGyhdxYWS4bPdl8JGS9tVrqJ1rp0cDxCAF6OvPgWIikce9QcLjVPT2T
p4y4AB/x64MBPFIfgpBXPmJjk7wgNZp4kzQUmhEgD4biIOdsw8herf4FQTMUUfHq4bp3LhEkZte/
QoDeMxeXH0AIOgnoErwrj7T35B92kFds5TZCl9byBdzutJ4q1KM4+TK3VRAOz7z0fvGK9iNjHzRq
/FXXmM+I5gNUZZujnEMNrNz3n1YMb1N7eL4EUGBLAvP8UuSaWPnQ+VjXyWVV7SxJJuAUqM6bUR2Z
vJFrwlduaQFO1tNjp8WgyxHjciqfJY7TsxtPgHT5TZTeC5VNe+sJKzYWJnLEEEOZHvPpkvK84xcl
ghj2gqEufdckfDb7NbDG5lBvCO8J0XRX33funpgWhoEhe/8+9a+w31wBMlSqXLsKoMxzJt2fk2au
OLJ8EOmSCu4qubolcb2QNUU0YThYHwPjR9zEG0BjUmWQFNDirM5WEc3kHmLd4mLd6XxvdS/GVfOE
aZLauXf/iWoFTn0eEV6k+OgbwP5PFG/SN41Hr8wLD6/tPkPosTU62snBir1iCy9sy57BW/kx36JD
0NeahfNmApDuAHS0CkMMeJ6/YhVIDu5ipYBjnosfGxilVr0U5TVbRVKxE8/aaOrSvRdmSUo9dWfq
gbD+Z15R2JJ9spccO7zXZPZtZFF37vhsEQFj61pgca6ut8ifd+H3V+kx/thoyBDm/hmngjsJmPwA
cicWU2u583R3kRLhpuhkrXJMYk+eXHbRhVdZqvIlQkcH8gJm0XHkpfpsuPn4EylEseIMkCiPmLA9
EBvKRjSh6TTh7iLPrh1kz4VBfVvvcaPCthZGuLcrbFvNCm9uftvFBHwlbYtpQjfRj/+aX0UBKpBB
d2TQaTTVxgkQyhSW+qnBggbhmurhjpWdWb5VfrpvX7G6IkmAUCPy4kiJ84+rRCCKij+4397LVjhg
qP4O6KqgYDZJ+MsPduzL35QjFp8nR0qXqtF33OSBMldGGCsXkeJw3dwXdroVicWOylhEMpdUQI3K
oG1cWFnA01/NEpHfFpsJRwWqDj2i/rNawZgMQs7pkdlXU3pcw+7c/C5BOqoUAxrDNkRMNLlWCyvt
ZLAWxIN1ATCYXGHVmF6mGc+6EODdClENKAySFKd9xuDGyFm0szSfxYkX6urVmqsKl+IU1CJdvMZz
CDHjKH/6Y5LjTZ4Y/IRmABlwL1+EyOCm6sCorvQufD/HkCEXwPc+JNWhnxwEfpjBY9gAwiVz2VBd
HvGNebYPPFDUPpWocEfd40swtzUMTgaPYdcVou+/mAVGLvNHeTcrWtfet75UeLCnCz2tnREKrxGN
SnwOcrdHyUaKzjHGiUhYA417BSDC53AFo7T6XvrZN5sxU13u4C2g7kAK6MlYPkKF4gGgLXPuhzNU
WQhGhX4ojMV2DETBGj7SFzi7r/ybUvzJsW0cQGAAA9jDSHFRU+Rt1qo2sOWTX4oOU4iu2Vzasn+4
mgAHtwJFPd3OYKX6bl0/3RBamvibjnipdP6kdDRZkYNzUmWl9ydjVBXdFHeO8aTxiMw1HurCDJGP
30QnIS7/NlILX8+9F9OnWUgnnq93as1jlFE3AV3Ti2ac12WAvZWmRJi3axU5B3sfH23xbRR7GFFj
J6cYmXMfdth3PZS4bcz1CPCJzn9bGZml/ZBuGL+U4QU5d7Q8pWwYHu2p3tIPrVkrCeuZJzazDFdf
8p47yvmFgrMnEvtVBfq/j5Sa29dGbpgNZv0rEJpeX2/WzE6RUfUlvrRrzxZb7QzdgT4JDF8uWKmE
sPlO32UjIQuuP07dfFQGh24HL2LnxW/GDaSIpvy6D/sp/pSambNfRbx1/Ht/wdPciFM0GHkjE25m
p2OnJhZIrp1TUVgGjKlX0JfLkVt5mfDLlpyn04EwuA+7Z6Jt9llvJwKC2ZJh1h1EN3IinM9CzCaR
pVhdHpw2xq/NaPKn5q0AOehGIB0B3bwNf6XoeQNx14HhwIXFC7wb9u1Rles+0ZvMACtyBl0uirbG
Xj6eGcwM/w6oOe+qdREazabxdKM/FO0Y5WJ7bdWr4swzphyn4NIbbH5ZEMRMagn9K8eB2UTPuwpr
rfPKm+6ViA9rUKFjfzBF+4NzomeW/KJvPfcsSQ8RG9sRu0E4O9XP2Scc3XSkWhCB2Hm/F26US8rh
xiY1gjUkfGQLxmJCXBX3E5rfqQwqN7iZ9fRqLCsPFLK1h56jbb+ue7wYtXS8C9ABhd7rsTcSG0pX
/j7AIwbzhy7q5juIe1mzEUetTYZOH9wO3SFNhuII8N93vT+cJb+ErtCILzaVkRvOruIzPegfqPDK
RPbNN3LhdaW8aBqYxr4AIUhASG3cA7tG0T7VIaY7OMtemkEOIaF2NEf0Ao2Z9NOMYHikihWTgVW0
knJShwlEC0Nw0keT5jwK5mkfGrvVMEYJgoNy6Xey4NcpJyHqGYgDCQXXhqxQ7lc3QhA+TVMspv30
zRk0ZlqEyy4Ed3zq7g3iSmC8hOTDnWKLJpkwwN2it1Znf1GqoiSy1h9PsCXk2eNJGwscjvSVkNnp
3DxKRWFruo1tEHtpLQi0DbBlnz27N8b1zizAdK95jkC17iOrhif3uubmP269Ftw2zsCG1QaSEuWE
wEGeBTUyY/MY/TPM8WtLszb3QFFSRXZ/TzSKQX/MV3GsfpIMJYxOIZ16VV4Vasl6Dn2z2CNMHWZQ
whZbbA30njAQePwULTnb+WOOw7n45RSk/Olj+iWJtXlLpf1RcEuyqCUc3aapWpfAHQQ2ZobUPabK
xBnKqJ63nmOPsDGO7fEZIPsSAJAbJmbwek+px18dK4oBfdIr2iATjBV0wodPI1nbS2C1/nrTOeA0
rz85l8KEBc2ZJedn5yN47TE1OPUE84rQtydW15uFvAnSlJlIuMQ4057bMHdyTW8vuFiB/gmuJaAd
gv65NsLJaVyS3/9EqBCbHvuIPP9qRpyFqKb+0tBXz8fxysWCpX9saypoMi5CQRwOKaRjFNVruJ/j
NSoI3IMeuFLK8kHrVDYzB3cIJTiKcPPDfJn/fYZkn6ZmY3PXKi3Rv7joXRBfHHBzeMW1GfEbx84Y
+NzysR59pTD37dhtf6S6G7wnpV8wChHdkOLQNOx1/8zjSNDnp/yi4Wtssa31yXLwhY/ek90kCBMJ
o8pD32i2omFaVSOfvocOoOtnTtzN0mL0jU3eheNHCLyWr/YQVM+LeHbWI+IkjorNvOZFlSJQFFXx
elljgrH3AwFR1n0HjQ4crI5T61wxisrA/wQmXADu1Oy+ETDXdpms1nKbYPJ/Dj0VskD4od8qSamb
DbsTjZSvFX2LzJ8HiM+kIG/uHZICv59OH+PDf8b42MkcAvqDyQXjsRxoZ0+Yc0qdj8bRlDTqaf5r
NS1/ufJWEMeT01v6cu+r6TV923EzzYmERG6wnOf6ToM8I8OHq3IqZujbwmiPoT3zDAaBKCE6cdZw
eRGiaPy9vovWFVYw6hhmIWA9XeP/YxZros0O5jbc/LCRU9ebuMtRZtkVSyVFyDtYdzJSbAh1h/sS
Y0g3XhSY7mB4Pm3e3ZtRuueKKDmcXUc5PPBFUGkAhl+r3kIf5PwMOEHKVQiYnJWZDokOHmppdigM
Ahk+kktemLSGf0zAu3Ab/Td1F5B18qwoBRiBSgZV0/Tx7M8gQvwJtWnjuoGYoDTj0Dk0kiNRjZbX
fkC5hvsZkiPEvgNilH8K9MhzS/dZvkZeG8cg3sqbvi0koe81gD5ag/cIOlklYD2ZXqAPdS+34819
EVuNKfu5WaVFjMM8LMPHXynyjiIS8NRPEnAqJXzhpnE2Q6lbLVAnUv2tycFInv8nMtxJ+8KIGd4t
qe8F41A3VbrASYjD78WO39cIYXZ1A9mL8WyUIJnfX4hlfmW3ysxth+gGDHPZkVri3yP1MmeVNwGg
ows98oREuCaZi0Qq3lQOX0SqRiHEfNAUun73/m1C4XB5rPRNG0/qd4AFXJIWLQU7cQbv2r6ipDsW
Nlv05Fy/2hlmv6j5ZEGdDGNUyR2ynftCcSKs6BmhhI8VVrLMe+ugBY9sHf6xyQWFJLPLl06bVBnX
0+dDd891aWeu2iix8hY2ht/GpC2qHbMQn1+s4M6DvQrL1TuTex2RTdSmcP9EYYjteT9cXyo/pIdT
r+ICL8G6Zckfn0qr0JIjrkB/i0wTWFa50poiSfxeSO5YdWEefhBVZ77RRVIAWDzMGU3UZ7mP+sGN
Xbl+vZev90Tb09Lzo8QVBIhQwgEjnQ3xkf0VM0Zs+H+apQaM0uIVRbAYg9babjSDlL7kSU4ivdvx
SAGw18AExT6G2E3qDBBjNnQx61OUSGNbYYJnp6KIE3pFHeGWz/TO3iBHJXJTBuPG0HvN+QskGJCF
WraC8m2yXFJyIg943KmjZsxkXVp9C8+90j4cbVB2mCLp+2X7omy/FEv1ZIlKQzh7+c4I5ThVLRAj
1uHpD2r07zx7tgBtaNb7+oYhifCJqKioSWLeB/02VmPEoKOo0d6OwjTATiii6cMAxO2m6bP2uzZV
Aho0eydK+H7+Z1Zqx2MdUAeAFAEiqyvuIOSEzKK98Bisj59FyRj0CoLVLvar9UvVs+K5pm1h0qdm
4ZjAcbS5BBSKZQXhcxhCuqbB206VfCAc3NYvT4RihNUOgn/tiyHB2ubvpDeTwPbR0nXMtQaksOtx
QYbrWdyMC7cBaMSjsJ+p8+g8dXlha1vutkRCpZ7Ssu8Ebrj/Hpg5sqKOWPSO6YpxAzJIX/DRufHP
FYp4GvgYPy/9/SysQjbCCQKdGLR/nQJgeCq+NSHeC3sqsIGxYu1/jtazHrXaqXskDhjV19XD4eMF
nrm3TASdtTw/aCqHwK5JO2kPqXFAL2zUPU9wYWBlgzIZ5Hoe2vaQbcc7mTahV21dai/k/MNiWs0y
1q7d+Im0Wes1l2n/NstIfoaTwjZ9TPl1w5nRc/2ooWPHMMyAt4YQWGp1pp7teYtCcdXf6wdUFrTu
EXAjlHJ0MMedDzp575of5dmwuh83Q0cgV1UtLSDZx7WpHZiLuoJJglSIzNwD1XXHLuBaxknjckAn
ubRiREA9r+B0UNkJS+vATxGq9Enm4vzPl1akmTK0uDLZHwgSN4scpkNzs7FQfhArWwCrZqxrknwh
lzjN8iQ5jeN8hsGyrS3NN1O9EVuSV3dNo5eddQ+zW13qR2E6zvhlxpuCa87+qny+c2kDg01Veds/
V6oCcxHdgIEZ5isUNN7/91Ms1Ya8H06t1DhSKGhqH3zn6U3SLHkpj8oxEmL1l0Qw/s+0F7C+F8nL
TXdUk/TJ98nelXaUUtfgC/l9Z+4yoG1Xjde36LGBeKUdFOoxbVWc99GWpl21l+tetP82G/r6VAsV
7l3RF1BDlMdDUnR0ilK6J0YR9swh0qhgZvHFrBeSNpmM/fcpQzLK1qe5GUklP1ihhSx26FuGynzq
ylKzuqUuPkKNk1LKuygtfz9VUaLOU3xQ5H3zPnqFd92ZIBZuAZ0UMyaXQZypd8jgJpFV+if3oyF8
SCfvucOMRYRLbU7kt0pAQ6lrsmKqbZDMXhwQgjxzotKwDfqw8J91gqXVW3nygAHfgmnxCfJG6ERW
y4us7gdlnOQwdttqxgfMs4dz7HqCNLxi1sNdo9x00f8b3etNOHHrfkV7M6MDJWg7Zj2N68wbhp+Y
d0YSj6B9jDNFqBSaPTUkZC/KDDJJzczmoJmrJ1oDwBarXALQhPXRIQk/zTh7Y1Gq/HlCc77rr+yT
3Q1rTjHpw1RIf6EghF1E47VxoxFf2jmm+tS0FPDjTt4lfLlnK6d0dgbT9RwdMrDZzhv8eqwA0t56
TkQS/nph4c38XjDH3hVTjk9UY1eFfrGqTzAvRGN12UHV1CJDhmuMum72SkOqr63AuLWNGNJR/5yU
RxcgflxyNeXU3UtGbAeXFXeV8B3LjIvMkkukN/VaCumR8S9rBnnE+52sn6aBMtQEi0XHDut2FmG/
qz4+QN+9qiGMVmW5JciPWhIVbqT4MiUJaPkMbRme0BwmaTjOAyeFvB4SD/fZX/Lh+S9g5GtYS3DG
VGvOtk/HQhIt0A4kP6qHY5jDAMtZbARvjQlY+59aANK/Vf6Up3srsJCmVh8BI1WcUg+1U3wcacI2
/Y5NaumFT7fyJDKkCWYbFXKI0fq8keDtPxWRhixsPTPNVYB/K85Nx0zCyvjzQlbKxDUvQOXcdsNV
BH5IW35eOWCfCm6TBAc19RNL9GXM+7H3wiW2VPjZ3vf7zF6WT3xLJ2/KQd4mj38tHI49hC37sD6v
1qu3KCRORLZF8MQ1PgB5p4MR0ViZwtCtMrwtnO5ZIXbSQTQE/zd8+sIrM1WvDSHk1wT2KxJtTPLC
3K64zcLPKFwgyEJ7EaxVKVY6z29eG6O5GMA37X/twRmJMznTIS00nRKPmJVvyZF5V6YGgrMr7LLL
kNr0laQDZh6BP55lCnjFvg7JbojNPPDwgcLGrQXNG6ujH+66vT9v2b7RB5dH8nrbdMGo0/MnVyn7
MTtE7fFsQJiqO/9WxyCwjGVrn6Re37h63Pt79iBCc3a8JlxtT83kCWBdCNaHoLhrc+HfGDnt1bNW
PQ6dRGlh7U9Ab4UKnHTodQcQJSyF5gPoZO9p26okWOFtbe8h2mexZeZd/RtM6WYPE8KkE+eIqa0e
ypRIl8+f0A7Wy3bSsX18OB3RWnmzZ2hTqkVpgwgOWIU83GMXxnFlDxri5E4tN9DWB/GRbNU/eb2a
Df7K2khF/QcbDqFl4RuLX5n2QhgyXuWWV67+4UcednHXlAjiSVpDtZvreuGCO0vIOxxZJ3f+Y6Om
Fs49Y7N3Dz1GXz7fMLyqaK9fjk6i0fW9s2ApW+aBJ0xyIiOQ/jlopSCdUl1rhlwT910lntGZ4M/W
Ly3Q1HnJpOBcU5kiNFAGeBtjaarcjckJYQ67LAfORs5WNPzUf1Hyr2y1dcCUwVVIL1GGIUpqhgek
9/ExrQl1HEC0NxYg/MrIM79anY3We3BncVruOMiMC3xCiHInjViulkXP4XhAWBcWmQhZt50sFsHb
VSK5WgK5gxhmqGIGwEZoc7MNoH4NY3A1NJpJoSX7A7u6RoKj3ZZy8APK1P4ALg6+WDLV0Itwtj3u
4KsK28OibMA35k2hNsyef+uK6HN3Jruu2yOSrdqT1RT44GnIf0/eJ/DiKAyl9Rv99e61yRI6BG+O
cqkb9kzANzIM72vBQ9MnHUhKXk+XcOjxEDWCK1pNkeKUUASThGsoN6HdYFpJ2+0na+qwwkAVEfQd
aSqYe+fT/oYZFUsCdZ0Ls2FTkfGqh4aM2SQDZP5ztpkP741j2wVj0FUV81AHp5PrbaePKp5H65+5
niXFWkl9mspzzIoB4UGc8b8nmM8Bm+6VOdjBFBkqU1jaXJ18cY8hRMUolJfcObWfmZ2VFQgOdKcX
r+uSksfOKN6uRdju34FkLwBDBUATBLV7iBCjJ5YMrbALo7Dp79o79HBYMGmTbZocZFdIqN10keQv
jpMwJncGrG2VGagfCVu8FJqjDe1gIuNg1d+NvodlhLSePUNPkc8VYORgzByFLv0pZmI7fXNp0Fbv
+rIQc9FqNiuv3TgPzKqajFME0Xna1+9BRJe+fEMs8dVnoRBMQ2hqlh3b/q8usLyPnoErQsxQePvx
x3P2gW8ct3IFlI4tLGNyUxsLcsqXDBUc+mr4Ca6P7vjc72pgo1FGZl6mWfaU5g/gET8DYnSUWgt+
04LUxzHw7IuLNTRd8manBQcrdSJwMDC0erdLkEo79XUQ8d9Lkaufv/AG5AeZAynQ9X4N5ayZWk7G
Hb1+2tc6a4LNW2MwhN1TmiSgPruA6uyW0PANCGppHAZ21DTfHOc/b1ShdvuPmdawmGAM6jcNcKfy
9b6CEurY76kfD2PeFmPWTh1UZXxFlpOu/JO+UQxYAZY1pBSr9v07wry4uC0BAA/wyVG+f5pxvvji
eC7AUHDU8G30YEKPmRl6vA9cL3ZVFIqEpyRSTsiEPX91dp+zJt5ex/7dJ3K4437EYyw6Xnku6WIH
+Kz2RjgRJnq2JXWGTmqWYMFllsugSH10vNFSgSxSy3bX5ezqVNVlOGc2WdG4kzCC7RSR8sBjTL1Q
9PTfKDRVnDNNCDpEwXviEm2n+SMRymetGXXMHSDdiarjnvRFuCZ5zHbwparIeRXh7FzAoiSn5Q5U
oe3Jydoui1JfrM7dR6+JpjvcV4tYzEM6dLk/tT2KTVDUQTqOfIKzpJSm34FavQPNxzLg8vkNpJpP
YMvYdNZSCMxfqLTr7vs/5m2LOKNMjoELHBMABMEb/OpM3HYsS1M33nnAj9hpGmMNPOClj0KQYEAu
44OETkBn360ofvKZ6CIKVGKagm5HEPapMkyinaEFiGew7Rcj/tINlkZtC6twaE2u4/gFs3rSaFf2
s0nO3iRtDwPTQzQgY5ApriZSNC17kwxJoAgzai6A/bzKtDLyD3IlzcRyGWa/n1RYi/qg5RkHitd6
B3fmWGsZi+LLvy0pSR3YoHAF9BpW/F50xOEgu71be59SV3jwd8hMv5aR1yRvaB2YJ+k82hSlfbj8
ELTGgeEXBDDVIUwuEBh7m5xay6WH5HMRSELM9J0AMPrixib9sZTCi6unhkC/wP5gMRrQXeMLNdZw
6JSSIpxKAeW06orp+BkouQMHOVQ8BivRRnUm6ff4ktllC1J9WdGZ2z9YhjlF41gSC5ayHIc2tiMC
IELc6HArvRrarN76pBey2p+YQFyL1yNSCbcASTIrOHQnWjND7RE9NYWzM87ugcQFPUTjFFDKYFMi
LqWpFJ8pN8Mo8iZlRuNZdST9yK8p0gSTM4mAzCS/gOwIJorOr1ft+epYRx+YUoEoxWfTVA9CP5dZ
rMcYNQPy/QPE8KsyV6jA02x/EFcpVHK2U5SAqhtRrpFuP1OLKlqzREwEUxg5yL1D+cdIBTQr2Yuz
30R5YhA6mMxH4/jSCsekpXSZEmyIjcYimjxY93fhANftAAkVAOifopiLZy/9vYQZ/wt+LIlODNoN
fYDjYVfHc2b/BwKQ1aIFgKQs+zJLjHoG7Efc4W7YTtTZBZYhHzcW+Ii585QbM3+ciT0av13y71j3
I/9iEJ8w2+X9IhEuZZb1KPpylmvkMoUbPw26EHJxtFkArUCTZUXBrYk6EnKMbA4mykGh/YLYFu73
/cr/TL0lj1vaq8AuhO8AmhEbYXhL4ZZpYCcoxD1xpIN8fn1C9jTPmZbHfNOM8K4flqGGAMVHqtBB
b8Denk8ZXuxiKBqD6INpLOU3+RjJAoaBUtzHgU8Lf41cI7HMowYVC5kNYnAbAMV37UhxqCZTzaQE
rov054oo5GxsA5+LMdo+sanUbHtbH2D00aTTqF/z+cpzyld45m7YO5q6Q8sJDg4IVSnUZ74sOGUe
ZsB4VJmhIFvI/IIKrLlsQc4zBVtUivu0f0YJ542rsD6V6wrfURZZhojAtZZAspRhJS56yhT5cson
4zDnP8XJk+Wzvgmxd0/wmcvwQZ4nv/C9Fw5lRntLPBkSIKJutceyYNw8ZqNTm+HbRhD4gg+FMSnV
alajvsNR9aIbCHdL0W+dqye29gMi+2ySQ5ed/A1bX20vxLTJSCNLSaOkr8PwcxPuTYk+s1Wg2Ghw
oEb/NicRt1JsaRIgffzUSKTao+pGq/ZQwy98lVO91knZL5i7wB9BCNydlQulg50WI5lB3wafOtaM
Ufby9q4dUyxXAEze0Nqwy+L8hyPqy3EKa1d0vklr21fRFJsF7HOH3ez+8BL1BXRLudgaS8llGqJi
fd6rEPVntTUbrrJstk1zZpxqqECxKg8C92vwOICMW9axmeF6DKJwrKTyJuHraNBHjOk1ibbV2Pfc
k43i6exyekI4pdJGw9CU91drIB+tKXTB/S6pOeg41TrAvCX78ypdmtA3fTp1bFb+vHAbyGQk2obx
GJBk4tjQUMsXDuXJqzuHl5CLK+a0SLwqFwCX0CsmTERJjt9mQpGDXw44ddjWUKNYFwzY6Q++j097
ujzK/e8i52tTXhxxWvoBYQEkXQAZ1dii78uqFYZHXUVsEhwybw2qPBvcd3qH9jQ7JF19J9+r/srg
An91ShCJAdvfvqkKapeDEAuOST/UpP0rC/hutGLpRGImvcd+6lEyqUJi79DBp78/EtFWS2mlRB6O
FOoqvR1J1smkj1TOmS21rDXIbYwcBfNuyE//FYER63CuQXwXGlPzkHkMdLTJc6pEsJNXirMR7Kfx
D46CXdS2WYXhRP6cakqKnp0KEBUJudZAirERMtF3wrwETDiYdHkZurkNczp1X4H3lkZngmgGjHs6
fKXZwofDOhuA52YiD+0F6QJ1jjRoJGZhxPoptDYW4DkjRT9DKPcypWL217X8EyuiqKw0wkXPt+0L
AvatAUc61cAjAKyEa80UTLkzJJctih9UcQVV25AV+2HaRVSo5aeap1NxYvIFnDgE51xcMBB2JUkj
KKB+SSOx526GoPdd3KHW/XOXjgtBUXxLtBxnKBIKZBbTdnOZsiVvZlA0Gr0PGbVs91BrcIjJOXlK
d9AH7PR1fph1pVvyPzIExJR1go0ko0HQQhHcX92ehxdDXI0dnJbW13jnXhvPYk4r4RSZcFo4nQrc
YQryDSQt5LesOh4ikN3voKUj/KoYlffG216nb2KNf6FcyxRZxiZ8lWouW1+cfcjtrzCmhk6ZBgZQ
ZZ7gcEceC+MhJSZf1yRK6O9GUxlOj6idtJC+/hYkMf0cmBbSeDTwX38nVzHJV/8yHUhW0OmUOewV
UgrgcEt7F3dzSfOUY5NL7jOqu7g3ZIBX3xkQcgcvyU3f3lrAGfcTwNf43s5Qt5nzn7yaESd+81Ge
DyHbL6fwkFAG+XxrdQhorF9BGngRCL+yx2xHzJvR60lpGkQOqJ9+6g0iJ26R8RAdaOoXfd/o7bZo
71DUbapwQ7tWAOESotmolaEBXmkk0EUe6e77hXvKkc37sXMOi722mNLL2207F4Me0m3bpGM5E4P3
VfX7trL70JMPygdoWwZefWwGImV20hIgIXVJI2MUxvLEpDJnBhb81e+2ySJV1Ch/zA1tsFGSIS61
2eG28j9P5xtMiwNx+2687O2ZT9pJNTyVArBh5pDVnxMuOU+3kkVp3R03zyuL6FTuPTFwQ2cgQYuC
//B2ej8vcajJoI+cVCivyd7yDdSgTLbW25JZzGxuJiy5sDw/QzS9N42V5cgFJkn2nis4uqQkJKCf
eb7vskSD7rVanKkwUuNG7ydp+hVGgyVyCXPGXyj2aOhuWMYUaeg+HQUze0aDLoYYks7K2i2tsg6p
HPVTLGDJSfU1/OXnYielMI47J6/cPyTRNiZSZLghDDk/NBnoNVg7VNP4rabmInXPpV/b7LikQNU2
Fhb7jN5gUxmo6y8a+jRZvRoAVv4kKqT0+p/PYUvyNAEXIJEbSCpW4vDdCyEVoV6Yi7RCVqcFVxwZ
dsj++lv3NNYhBtMh+8YvuFfHlmmKiiEJA8x+2NdEC56YcU9MevNOh4mSdBQphihFlpQwn6Z1f5GD
NFj0cg6z1VqiQBMZmW7Da0PXXD7ecbFrfEAxg2Nn9BdgAqFi7HuUaQAbhaYIGWtaSLo5YsgQXesZ
nMh3zrjbJvuONluXUtKlb/e2HdD+uYFqKt/Vh0Ypc+xEVxIbwFNCnpKN1f3UomwO1YEzz5d9qWXi
/djepMFvc48ADIO+f7JkHfV4k9Nsad5CEDQdv/a/rZxeGsIPRwPPKMQdrzNVzN5UGFVfv0A/fJOc
qSmOhyJxNS3sn0Na883oXxny/lvcyfLHX1B57dkSBd/NH9Z5wpe+G2dAvxtFuz72TzhVxwdmkWvN
KoM1Xck32Mobsbk4rpMxyB3EeoX0wyqWIWCB4BRKkwfjZnIh9aphe0avGB0szUMAYRbvNXiCFDOM
BRmdImog5Fyk7qQu99RXLJOMGDCxGGQLeLarXHBVuzULMghVB0L/xo86rxcOy+q3MqrqPH5MfrWD
Bca7oth6W+MPdBhnZldQQHH0bD/vIysJdx5vXShoni5XVC1D+HPhdcy8aPQZdVZKaxMGANZ92Y+s
jzKA40wKSneE7V44oz5eyWTtmIfyw7TkR9dWrtLd88B6hp6GN+iJDvH3v9C4EhO5HyCUFK6FgViZ
8Nl0OHkV54VNC+3fB0a/GFgqU6DZLdbGqTuapJbvRhinw+lxcu00J8VC+23QMsi9GlJmsBQmy9rL
NTPQmwPyKFTl+N+4dNZCcpbFC/PI/yLBSzyb2mwk94SawbVfdQg9xbts5GMuY+Vucb0VcZ1em/0k
oSqQqFDHIhfcuN4z2IecGK2Nv5CX5R6KLbNgbu0PXF40C1CzqsuaorcG5nDTg2ZiqJWp/WjEyKz2
2lxhD8q0b+mJydOcLGbj4bbXgADlCXwz6OUrRAw+a+ROw8+acGBhjGULZB8al7CT32G/zQ0+BWsu
2vREzYLnYadxbSdZ7mDQcefOT+AAL94erGyO5X9XSdp2sZliww7TOvjlKA5Gi5ByrswjtfHZdjOZ
BRV+QmVUyp2PzyrWu1v2lXlkaT+MWuS/HfsK3uN/1ZKjBm8NinW444ia0iWKUWtRLUfNWtzLEA4P
6C6S1z0lAdVGftFs3X2FU0HI3SAKGSfj1kROAIQwXHx8APugrlh1L/atOAb9h8HiAMADuS8SNwcf
ahj3CgXRsQkPt5sP88XVp6yX0pJsnvVONUMogOzWTFFRYaQ8W/LUtgqwvFmFlCErbqyGK9Eto+Ej
VUwHc7GRUAyoYsNjfyRnNO5Ffzmv/qvADbZOzUq8fu/qC9qtRswySCDR/PYKGebL0Ix5tbkzXnxH
2yQHTjZKNuo3uwpcptLkIkf4KIwN3SpYqW3kfsdlmJik5xOUYzgc0mnXqJa6JTcdsOaPVgKga6Vz
h5ug7WanGn/G5VnB2bi/GOZ9D0P2B+uALpbcrKUPP5jO5du9asu0Z2EzgumnUB8AYsBIeq7YtJf+
icY+Ov1qLyzZNrULsdRKE7safj/z8nxYPJxiA2SgvAhBhMwZJQQqpFEx5zhRDvV4FkoDgJsaMKZ9
QMNrPH3j/lpA0q3nhN/0MRa4lAHvScK7lcXG6o9u6ElLSAjEfd0DDdzoW5qvrx9RXEGkVDxSLd3I
DoqXZwKZHCT/J7V/FN5JS/t08icPJql8NTn28gYpn50gMcVvGuB1ZUZpd3nKILx4B6SzSb5ef5Yr
cPKLLhsXZVdKzsnmuCQ7JLD+iDwm2m11f6lDt/eiSlkv81WEJXFKiGGv2hwK7uCnVX5VV6Mqa0s+
iyACPo9V10iw2yKcvcVBEwTvr21ko3xIgTgSbmpJBBWAUeulVGmpENsdrEkD4Rt5XXzh7eQG3diu
wO49z9px8F8vYWiX7D8AJbW+vO7kxm8M4i27+b618BuuLNpPquf5l6Q7wjmzJchIEBcfmI6MkXWW
ROUs28ocbFh95MGHuugfhToiP7h2DkSRLwd4qAxgB3Td6X00Q1ZdDthnw1ylUVr0NOah8hvQg2yT
YtSyFcHOgB9P74XDIjU+6/KySXQnYZ2hCAkBLAxK3rrBsxkMAc5pPwzUd8NEv0SUZ3DoSdtHH3QJ
SUnBuwPSN/hzDpfyTTrt8KEqggi8iU7dtRIlK3Sr/f8Cs/wbJoklKXTgj/0gCRjfb987qfWta67I
cqMmALDIdbHWncnavc7NvJzcdJZkbKx7xY8ytHfpe7S5NaELkDMKKxTl9yt1CYjlNjAIkklgM7ly
JoMcWroxPHQkXdVSPuX9O3w9xDToesEnAdLSyELbGYWB9N8s9eylEZ5M/BbPZo7t5Ft1gH9HWML2
gnMnigy7J7ADe7gEn0yyJHWB0CohXJa1znUzYITbzxXzoDFX8dqgZ1xObDOrVFe43AvlLt9nWvXC
L7dWvE1pQ/9bgSjfcNrI9/0RtcUbke6us0Ij9pAF3kHJPjGBt4Tqjo6QnsIQN2aDo/L+Y6wWYp8l
S131uYpxbm6NNFRcVIDOO6F56pl5eOFHiStSOCJXL1IRaR9OIQBPhtfBRqr0YxmX4k+SbeRhXxnC
8kbXDeDavtFCLY3j2rGOEjcr8+hX+8wTwMwX2hSlAr5OfLrWxTwxtPMEXHN5ilqdFl/QWyt3QR7A
bufEQPjhH+uIZx4xHZv/swr2MDT4nZQztcsGg6MeW1zj55Bp90/Xz7JlwuBgNcjjw8JNoWL6AwdK
8yk3aul2tO+foX4JTD/s+c6dS9Ua6vYjxkaqaFL7UjjQBp73SH1grSYUohgBwg7QR4nryI6i6LxH
uBz5TUPXRb05fTnvj+uhBhqZuY5sewsuyJ/Vp2tB+wZueboGrA6RBPRU9c0ssBl09R4lkgXIzBba
pKmYRawjqsWejAPnDMxNLLP2jGh3rjqh9wqt/CZ/wsxeWdMNUJKZ9PvN+wRRhmgPGMUO7eAsqyCu
oHBTmlkD+pt8E6e5v3GzBVjzhDSu382X3jrKB+3mgusDTJLoRm2BcLaBRQqDHdGgoK0WWc/mRQS2
SJIB3UN+HSVOmZCeeK1TwIendClN2sE+IAmRXlvIqeXA7c6E47oAfIADANpK0yCt0pvrVEKHvhAS
GIwIotKxt0/m2DK6tKG22+lBTXdZiPD4uPC9e0MpV68V53QYCSNPE2mvg+ndjPyMtmfg/iptvlQR
5zbL1gbhbZsXx6ltFm0lKlRoFBSxarxDHy1XWnHRxyS1Nq0P2CRcuHug10TFkuup3bRN6rkC5QvS
VKA9wrvWqHx4vS+zCU6hukMWdj2WLzjbTapkLv6QJ4iM+3QXvLYr8EuomftXKliuKAdGwRAYH0Do
yRjZ0rqhCu9nkivhIIhQQlF9/Xe6llkLrJWvmwEgGlF5I0Lqdsissj/3C9CVR/q3DnvZsJFLP6uP
B1NZek7/9+9ytABqX89DGe4AA6oPV2I+zcgkjTE7IXXO/8mqNdRquDP0HSdiVgDBAq3MFy9Wlqo5
S3z+K0zy9rohwx/chiUeEgczl+TqzPCozc11pNEfYxaq6UE62JpVjCTdYghbEZuJAErYOb0+mGTU
FHR163sibhi+1fu3vxzraxDVeL4bBTiTYXrEtPO3zmLjf1/bAEF8uPK8lAWgZhk+MHaAW/KOTyLv
OtYOZ/g/xi1rvO7y7HBKPUqLmPEuhwGdJ+V6MclKCTdiPygQxTORI9+l6ZPTMgalMzEk1VjUUMIO
gmQz/KDymFMkPmt0hugUCfrEEQmwVMHO1qNk8Oqi4CmNsWXLvgyFlcmWZ19uEqOxzt8dvGCvHPZh
wMhtHWWI6zLx6o5kZrcnK5m5RcSh+/Vj369zd5vg5MVM49XmkRMDM1Ee8SL58BM98vLOv+d18oxH
81Pvl4BTM3hrgi1claiRJx1/ZC6/qR/6q0etRhTg2BNGA+0fhHq8zBdAYfAI0XCoq62WvPNtZRSn
2jHvCAxqA3nWx6/cgkhOvwyStbEP5rgEAz2wRKpW7zb3JWdG+PwtknHO50v3xruILBtkcCPxo4Y2
jz1sKQLErig5y7Ep2O8vn/gYm9db/fvjFdKB37/n3uSm0Zl4POQeUlTSUunojXh6MKTmTfbaaNEG
XW4TIYdtv+cKcfNTiNR85UPZ5K9rarlLLHSNpfeffeDnGYsAi5B34QB+X8RSDUQisSGtNXYp5cpI
QIXslq9S5A318ot8MzEDOxFJNZIJyTCk1l6NCot5+TlxX62A0VdmJh+GyPulUKCrmRNKQWmbeJfR
p7z+uaxIOBxGVB2j/iWn6r2qkbaTXtvb9Cpnqe2loFvpnjaLczRAgZxq4YhgL5sTZ6uhk6QDpodx
Ax/tgMecV1Q60+5rCMIR9NI4HS8miqI+sCVYC5It7RxrVEEN7dl8acfKD2vwD85q0IcR21KNEpiJ
kBtWi3AVfYa7nxRHGHq4iESsW3DlpS8E1gSCELYO5WFSOEzCnyYmss94IGnAVJVwdiDioYFv1WFk
AXftpFMnY4Dpi3GNAJ8iKos1PhEtMkqHdU1OW3CNXgA2KPkMy3Dm+lNjpHe4fjko2LAzqeP8QQ7N
cN+2045BT+3t5haaRTfbmGRK1lCgta2HTCyBDam/z556GQll+aJBoX5koK2iNyiuad/M0gbGOJIH
IgikBacu++dba+EbJhyflqkjROfKl4JRZfFFq0KfnslWd1AYSxyx4jAzUMqHpi7nNfZ0MWAP24IS
WgSCUuwq8gHn3e4hdTIwzg9z3SxOXT24Q/IMgsfP9eF3zB8TK+XS81OCAMMV2s1sy0WGBBKSiE68
vUMd/usY5yk9z6QC4GHpVQvWy/IlTMGtFjITEB9/SI8oYfYktDIcyKSQEifwIMHvN5eCuSCoC/CJ
yA5zTghuiq3zEzvSzkIMeAeU/lTwI77/VipfuniEQC8LH1H8Wzgj8tKstigeCqgRngqPtpoO2pUR
8jT4jF4Jue6bprLrJT7hK7Q16im8PxcP5KL9tc8d4fI0mPJ/tu9htPDDnPUGpwH/UzcmnVk1OJXJ
omBFdVwqfRAx0SoNblwwzqWFB6AL7R/+6HK7xPmPKq4wtJZXvqbHpX/CsdiCoGGjXxeZkbeBSg14
zhhN+LdpYSvgsGaXRr8idTSeB1KDpASKQvrL+ufRYdY00up2VLjrnFDBhcapF1nuKOZmy/bBxcTs
v/iPeeRHJt1R/+YQGp1bQwvSpdkRfgPwnlSMYxb2e6fw6SPRTwPf7kBTPvbHJrfApFZ0MA4NsQOa
26n/ycQBoNlJGKK4+X2tgRaNrpQExRz9aCQX55j5N4qTFOw4bBnNQo2Cjdw3pVQOpujs+3GkorLa
qeEiJfIv/oO25Wb9l1byFeY+f5qdOI87DtVD5RpgRIRdrvn5cG9bQ14w6FA14rwM4el200diXfyM
L+tnIJgRqzHjKvVNpeSQtBJlY09hFQQy0yjlWwqomk93R2MdjdBLuIHR2UweFaxBBcRkGfDxz6PM
09jeM52sX/Z3n695ed+AavCQ+1Kr1DbIYwHlcMu+j76ewbnsAZ8iVAKG4alU1hbc2X4EA8FO3qvn
78woGKGeJqVOszBYfL+HzqnOdfB3oG0IefBRfOfMitW+nBQQea91FyLUg3MPx6NQ31lHQ4LvMiG7
40UrNs6hQAIgj6GrDy5wX/coDkHTslIG3+zOpVEP+D6R9JYNeokcaq0IIGDhPwyXblTW/3ca+I8X
zi409aVv4eF3GjLOxUbEH6Iqc04JvMi29eOaP/8sQ9wa18jvr0xHMfudciLL6mmrDXWuJA2NuHKN
6Swjz/Jsh6T6I88x/ziTop8KYCc7qCSBrUJVR/kGPXynkN296rmNM26od2b+5hAM17yaUWpbcGQX
z9UB709Qp+Lwm9fAZ4IOvummKc1hVCXTuU8+iTsmDDl78ella9pYl82dRqF5yZinCoaUXmD7MQJg
BCTG55VP0v2rTK/NAlbH8czl5Q6kAaM6t+z4EuF1vQoJO8o2NI+NH+NTVFe9jXvmive7SNK5KsB5
fusE4N6ZUfTww5pAFOyDOMJmxeE1v8iqT0JWmziJNnIVE1erpdA0B+57n1gg8fJQbrR1YMrQ34mb
/kxd/YQacbpr74RVW67zdZ+MmpMsbkhidhvF81OksKgDEyJYpEIFtOIywsNGNOY6OgFdCGjgVNLx
/3wHdVMIrtGUfrIfSUUGDR0VG7cEOa3acVqjfWxYDurPgUxZ/wM/JCu2jLzN5PpsmGMz9/R/ygTa
CMty0jsMDlPDwEs3AZb/qIhrLls2CVFroTBg4xI0z8MfMpmJgywqfipF93ANuWgr79S8b/mvxn7X
Hia8/+9bG1KA7KhgO0b4W3GafG/LD70VWvl4s/iIpd+Spy14vj/SRVpG3AtYNTXQaB3ry2uVa4cJ
aDen9xH+YLpjta4O0noX8k+Pt7m95eVz1yvB6uJxyD601xqx1uhXx8YMnrUhaADHqC13g9F8NYEV
v48VwrvPPimP6V0jUKK3+Ob1XqFygBgM/TEsmPKiTGphUS1W27CzKZjSLTWYExnTnnWyPxx7Hazi
JlZNMUI/qhKEkMFptAjp46chEuzPtJx+0ibaAdccBtY1gxqg1aP0jiKk7Mm1Pxg/0qXVnm7jbqWn
QvmDfsp/vCy3TjtHVAl954t8Qza1eKBGg4PhfsgmncC4+zG6zLlHz6UGzlDXSUBA/0trMaLtSVLy
hBYUJv3DZ8puQdP5K7GB2/vhmw3mbZEP5OAjucDc60bIpAaMN4F4109gPJjl1Sp5uzDWX6uqwMW6
tqA0/c+uZRsh1hl8+sIVtqsNiieNEBQdYl/cMHtcwngI555kJbh/v73xwh3w4gH6oifQwlVDdHar
LnG/leRNEFhmk1BkPqPbTr2bR8wApJDscw8OTl7jbZ31SL37hjR0qDOyZc4EawcORHKoD5jHL/GT
kLNhnz25ZSjqSOmjcTlof0LuiW4zHNmewjdxLjac2WXdF5JeDev/036Z2FuFqrKvk9IugbjtnJx5
qQGgjfZmMXuxmwbqhgCK8qaZy4O+SklXknFeyaTcC2E0a4PXdjlNsbzhX+GxGsApfRQ9gtJIeR8P
Gln9WVBZFPGktptQWRfqAKx3Q9pqD8PkGggkhzJkRgixwDM68ibWQ3be4vdkAlj8TcA4LeXYeK1I
XhRsfW1Ha4FPKuaa+ujrHFgxWvj16IneKifohvihMyS90W9/rk79mSLkEI9plszRCQwDzRGMJqhP
aNfESJmU4Xe+dPw3FhaefxDNgK7GW0FHIeNu0Xk5kjRtdqUC4s4aLDyXXwIzbgrl1iNb0ihimQeu
CM3i+WlbEnMDI0liNDACpziAziM+kjZ9gh0sfY6ecubD3OS7wKUqBzfQqFcUR2+Rj92Nya/bUKPI
SfHONeVUOZ2ePSrG11Va75uWoLss1xqXGaWvkwkMEnsTuoY+pv14yiquwRyRzYc4fGwjZTniJ9zy
Y08frAr4UCJ9UC1sc/dfkvCX7pKDJRPs5LScmsGK8FifZ/PY+A8hGSWKutjXrAs8U/lJswPNCUGY
RZf1305yaR0jyFa/iuL8f2TDBhzmn4hSUHGJqWtrsHcaxIpPj/uc7+hA+lCj0VJDOSnrjbdZxH7X
5PCjBjRcaNibMYSQlWfzfg6eCVqjBoxSh1E//l/eN7oN2HOW+8sz+hK0DiA8IN82VlE6F+Z55/P9
Pp6bBfXBaCJtlM5yvwbofFa1kOrIi5L04Sg0ZF6RI6JS05VR58BoJXBtVebT3iVuxKl57TrXalQj
N39d/9ZtD/baZFTya2qjOs4zri8LTlu/lZihh/wOuqa9oimm2RsKuHwdSeco9v1ZIeR5tgWbFIdB
IoxgL70Hs5E9hupMdtCs0+fehpTQv+WbW9tUHLYVexJ3nkuelkvmritZdZdS3m63/n5L00x//3sA
7N6pyJ1TLAUtYESINjSET7VM9t8m7vrZk12uJ4hjoImKBA4PmP4riHL2kYOA6anb9paGLnIK4f1X
+oEdsKHMJoqM8NCQ1RkEWdgPxAfIICxNsP69sCE6pDc7x03mtNBv0q/Vb64vrA06PDtQ5fhmrHEH
Bdaq2SZ9twzJKjmT5uYmVzBAxy7Y96RiY0GfxAdCRTsWTG+5CJrwVYdH0W6TzuugOWnUrVWVHRqg
vEtMTFwV5q6FkJWhvu+KduWj0+i2sMsX9ttnzqtENccq931MT0TAOh6LkgKF8ZB1kc5R5OJgOp+C
a5PDthCZ3ggsSK8IzpY7EbmJqC85Y6YA5O8dy7doeD+HDGrBWQZob4IU60JLbZ7ZfkP974zq6eQA
9NWd/x7Htke9UFBPRRTS9HsUSnhN7AZ853pD8aXKZ/Zg+2aDpYjP1bNX8c8iCxylH2/1tWAsVpym
XNzRR/hb7p2uGBJv/rq/16fbCWBjDtnsRN8WclYmDvwGg4e/2EvKaaCVgYWeixaCjqStt2f44Lb1
KoX5vhdPSU7sDazYpXXUAIksRmdEHuU0rTGexuIjcyM//HsXO355xEBMXFQNsRUnXGG3wjQA/jRL
NmYwpmWfk6JFIeENn7My+H8IOQ4n/tXJP8mDvwxKYY7fobMx06Tn8hN5LGwI3jDfQ2+p1MDo+FZv
EHzMzB+HSYP0OypXjrmRHSUqji8A7DJpNfCfPE+/802NgAx6OFf4VT1hGz4yGDHRh2Xmq2yj4hz1
xAbrvGYb+RV1oalVhbl953jdoNGDodnwAzX58qJ3QbDLdRD5iX4bnjI+u1wuA0FicvSpf4/9PtPH
We4WCjeai4PfS1cH6mlqinJvzJIOGDb8H+BmhEGbE/hRLlvesIRWCfs8shuLxjne5q2bN/Cy+J3J
B+Na2DX10t1ki6eITsjilrzq6P0hnV3G2+b5nf56hU54iepRWcR6qeBtJqNicnGD5E7q3Uxdnfrr
i9cUi0cf6g7uyD2GsIMMtR4Rc1OWycC4tJEvyhI/7lPNDndOK8wBgVU2UH86SENMZ699B81cjQ2L
pEb2CSPq/h3ZlbxRUZ5QONvYliawRrNrd/++dp8ZbAqBGcaW2mHz9EOk5Ani7D8cYGphMotbmNCg
twnT8KkxrJYQbjLhK9ECqJXKEyrUGXBf7xr+rQ6HKMpSJFbzRxtX7VvSxKdYEzJSguDf1SzYllLP
K+KFQHrH52MyRloXniuLr65E74LCpI1bDcAuEPrUtQhgHJpf8hWhZXPjYG//WkdiYw1mSdOAmfWE
dFblwx7uZinXFf62S7ta9HG7UrKL//3XmOrInaCXzRcGPmFQb05N9oUHmOTTo0E/EEfkAJiL4k9w
10jWPW0gEdAGYVwma690lMvMDxrQH7s5kCKz4ZzcJ9vveEowE59CL8hJ1VHBfaA2RA3vcbWHDRXA
qW/jI8/TLXg6tn3Dciwu4RM4BfbfiSo1ecBSSu7r3TG6gEROCxOnGUBQwB/82+zQBtsI+zMOeUqS
wVNSstQtyINxfj1h5z9R23uDn8ax6YObdg2s6k5hW+XkhLxLCMciAa7zuJNFEVZmus0jIylAGTFk
yULBmHywBHY8gK28uJhvfj+MZ0uvUIlIWWztF4Olkw+4m8CN7MjaDbNDOguDAUL9JcGCsH/oTwUg
sdwEN3GQAtmNUpXs2V6sj/hIEECm6EFFjTlll6sRvYDjRCwnsu6g7eAeGkRDWjmnmGbymI/UDej6
++6iu5/QxRSAam28eHuDySetSyPvtRyQ28/xMZEPNaHDp74qy0mdpyVC45okK3bWzW8MJ83WtGAB
y9si4VEVUgw4Vh/saZtbrLtB1LQbnc6cWVpF2wOceVaYzGG1iusRtVqOmawMmlagivd+nWArudug
cfHB1+Mj1xeXSuKC1AReSbuAAOTkt/bUUQcmudVZcIXp35hc+Dk1kzXbCpgoOxJXODaR9vkNoIIq
/7OadhBjX4A7l7rT1dHdD8WDGpfdB6szMIcimB4t6O9p7WtOXga2U6iIoEXbMQxzgVInWxbnwHHc
psKeCU7vZL9nb94al3+IpXRXmi7eAx0dcabdw5ZlJM1ePGFCs6SrORwCev1GxoqlJg+voMjB2HNB
b1D2/2PbWwfjJw8HiGCAaknqVwATAo4REyXham3x7tipWvqKpxBJa0DnCseTyTidPLX9ng0KNcKX
53m+BWrJuAX8guCq/vSi5VHaLNuZagE3hacC+Sa1wASpBiP2N9yrfFoBtlmS6DTSbUKbE7aZWh2b
W4XfZMmrzbu80j1lz3TpBy+3r0of4lLxf4hKcHQPAgKkWpLfq5uyolJT5ojLDw6w91h7tikvPPBW
kQcvoZtay7EjwryJENU/zRVN7CMoZktZ48Ef6LXhC5CrxMjf46y+rUn8zmC1+mvnGPy1C/58zb9O
bVNH4ks+lXP629/Bt4u8rkLpdFQV4q31+10ld512QwBgUF6Elt4qwYWw++Im7cwxb1BGSNEpxxky
F64sCvXSLyaTGlEnpe+C8r5UpHvBfQa0qyuANvUdUYfeVfoTrkDoJy8Kv5plOD4nCZ0H+R1LM+ob
SKj8ttfEDx5soZJ7OKA9a+X/dR0ODP9YKuqIbUt0d7m7LnSjw5UwWV2+h79lYE9tidrbQa1OY21P
HU6nQS6nI/QUlnOWnKd0qVa/ep2GH/8LjI07neyVfCJh42LQMazTLzDrjRwZn9tuozw3kBEZhtTh
77US60pbLF9Ih+5QfnOitxgGosDUhBa7DgjgXaa4HrmUaxU33BaR8NSr21gyVtz6anE8ihVa3Epu
bTI1mt9Dxn+cegqSPdt0LY8H+pGd5kZ9T9Lp0pYAi1O2jF8QbaZBqH2x8hJdPuLeOouNYWCTBuXL
6lzVr6bRiNoThxevfViWRTGWcwz57YQokddBlwyP3M2gk/bFwjFQ+q5jLVs0hRG1Du7O11wqYe6+
iByrbtVHVuqwPjePTWqGMKTuf/gbNXsS6h8T+TdulcVDW90oHysWWidHBpMBh9H7aKDrYk4isYYC
EMbI3p36rCqqplU7pAq5ncCta8KLAfYlnvO5gtIKZgHK6m4Nbr63wqD6VxFtT7eMvLt6FfJ1f2eZ
PP7Fl4B3qKNJQFEZDaY7MBcWXwabEKJRacBqb0KRNJr4iXWl3hBiHjGDElqsajn/VZfwiQymSprV
IBKQweFbM7Be3DDYXH/DOZ3xOi2SWy7aXpRsNw+KWGLgPwQrhKUdVX5YRXmNLFzAnG+hcZfj6/OR
7Z4ZLuiIdiL5Bz+au0f1X4X5ckT4aNUhCCvLFe+RqwCfiLWiSGJ4Fwvn7VJutmj12g7aChHL6oQ0
ZW1ZlJEY+qqSN/qTJhimVIS/btGPq2a1lOhSWyGgDHZyh2scD85IfrAMQT589Yk5oUqE2GSn5bIQ
OMCRcQ2AwNHWM5ZjjITxk7rFrvDIRdFafqCRgxQrdX2SJR1mIiUBY/u8xUHif2biCSwWvsvWG8af
CFFCp/NzYxuRZfwP+3zyyLww2N+MOHon73juxCIBonYmK073VeiiBf8HCqDpzej4ABYSpmEQ8Vyt
UR82+Mo4jL85Uh+4AbNPK6OE4pcIEN48UFpmpivNer4SnzAXzBeep4zL7L+FWPjAgBFKr6xczAAV
CMl4xVx5aLoczi3M9qrHMKoCWa8z8mauMCuQOYOUYpirmkT+31VHquCsJW9dJXTVVsvNElh0p10d
6gJGveYqfZUUyLBHfE3bjg7mV1ATbaCTwELGll71yokuT0CGGCOm0bGkd+WdcIUq8qa0uYr5kRLA
EwgMzzwIe+eNWGr1mrm3oZL3J0/DvuvmYzmVId9l1jDromZeQPNVOQ1ES8vCDPLM9DPBOcGnq/wj
aiJQBw6TMGaHMLsmULJid5RLK1+++/nVl76gQVtBpL+p6pWcaUFbVWToe50gRxmivFBkctELRVGx
AFgRjJ44hXV2ojnEIGSQfOb6xAudEw3aHH9CaT6UXtESbT7yHec6H8OUx+DpAyEFHKGW3I+excho
j7e5cf5laORJZ1zkfuKSmCI7j1MeW91YsOtoTfBGWGaBrcBYzI6RAPdM4P9GOZNbAE1b5OayEaKr
xZKtVSDHpStud9Z7r/PrphmsKgZXSGLP7RIX/IMKnZRPZKThOElnjzd0B6L0VZtd+ObNlldOyZDS
8e05Dpb0DodMd6kriAUy4pj7P1xwQXk4fitZEijnVTFQenOYARTaOcrgSyWJFDOXarGWsTG93BHj
jjyVbLQaiGlvom1FBZwo1nn/x254S6+6P3KCrnyeF2XQaHMCduQfXpgGgcmRviQXKOfzG1i0bkmL
MpCyWqI/E3VA0WYlwVi1dXUAOlsdNRv/sNnl/kJ7bDH7e+d0KrvWnX57nLqgUVDsEnBue9wNg80R
WeRhThUndsqoedi25YsensWvYrKc60g2RBwkhjvR+bfkskPRJqS4whX6LUxZoo/soZ1gYnV+KwIZ
F/1wFLgfaeCcqQQBlAAssij20Pczev9XnH3qK4mtCW35ChSS22lZrUIgUE0DaSym/DlwoEC4HY8L
V8RuOXLtoP+5GiYYJtyOpujeU/f4hbWJVsOOAhqC1cqAwmRLRXEyG8ycCbxcw5iUKvVkRdcf9kVd
dk4SKJwLK50iGNGlIb7S0VVIkzdNgxVOjj2QVMAO9gwabhpmpARI9ksE84SmFnd00GK1kV5wZQhS
gH0dt21I5/Q71B2Ssa1azyAwyw+2/ORQsHQBLErjIl936ZZONbsIua4yf4JDsmANrPxhNSLVQjaE
zEJNoMoXwMKD8okn5LV0HHKZnajlpjMMlkTnyUmkUiuhRpm+282J6OEVNEfagLnw+oCa7McBgCsG
4+j7Il0iUxJ17qUOcl3YIkieOlPxOVSqcPTIgvFA/Jp1qoGyTEM2a5YApOiVLnPY2Op7v5KvKsyH
JuGr1hLOBOvRW5hVUmpdhvdTqmLWxrVrdeS2N5YXltJ35FxyO1ywGP7haL7TKpY5uuwDujCKj0bt
WDSoPQMTFBd41W1XIplp9M2tTxe/9CMPNuJTaeF5YJ4wcbkk1XjBWqNqTo14LuWPwj49Das/dYiA
549TV6wf86L8seWBr2jlt9xwuELVyYqL1EEQAx15K+7N42p2zwz5H6rewOPX2jEv4GucKkkIoF4W
ZKiE6A8owTHPuKKDAYaZAQOL1IC3d5Hq2MtbVgjIr9GECATxjJZNNTEDVrA7ULJgUb2VA8zYNmeO
wTPOep0gV+yWnAGQu0CS04+RjLLLFrzzazYydur4++nY66oQc6/7iOfyHGSIvg/yjLFhqt/jChAs
FTAp/4nH+0R44pO/2AnSbrsFCBcSWmOl8lWXynOgGmHjOvcwkGHJdm3OvwHHFJ3hEbmaReOxG69X
27Q91/ermCgN2DP9yeV0VuLaX9D3F4vA0GjjkcYUCTKFeWrxjQICXi+tdsJULv4RauldTsi/718/
c6KiddcgnPL4WmJw81mPj+uDpBw9H1ommYe9ribwiKtTiF+ODVMy2V+6anwTSPOgaI5tVueTT+iI
3CSb7o7jGtHCJy+E/K7qoRKDWF5HcG+xdPJntJwd9XFAnDGB43ROD5BgsYrm5nCu8mdPiozGfZfx
BHY4uEGl7dYyqlceSL+6gnXPf1aGp83/H83GIvqtGq4MTGMqEfiXo01M4rH9vkR1orfPvwALf1SF
a5QBXq/LYDLaQHUyGnQSbS7oi+Wu5rsmmo0LSTuATwK3h7qRvr3nhTPo1iaM6sDXo0m6PKfDmrUm
PA7BKYhMPSXh5f6HtS7NXwY3huTx2hCLdUgCTbLiBUBZ8DQtt2MqLXvWu9Wp6Wn9AfnZNkFXfb+E
5BKRnble1ZGPHo6u5Mx6LCG/Atxdy5P0+XibTjxnv3ZWgmQNdXzvwSKP4dXPl//YZiBHkJPhzIQh
1HEg+omS3vCVAN36/+MfTAz80Oeb82vwN7iKgumGDpbHsPzxBHFjp1+T55jRLQ2iMwnQbMnPj6ch
VhIOJq8XhmPBkrAiMGg2zhVGazdJw92sKck52oO93e6ngei08bswAIOuhYcCvAzwBFoYlT6mklkj
zPAcakkSnnsRlnYrZkugWj/p+w5biPktVMbvVvivPqGZuKmIrWgIUPg98g3+JhJx7h27zQqlmf94
vL9YzQ3Zw3vAN50CAry0O0M5q8D6WLptHDFkw3Q3o/lENhmlK3gEtRMNxwTnB5OtZ56tStX0cfIj
r0xhFQpK3IvxD4aUyLPGHsSB1svOIO+b9H+GboBJGhe7z3E9gqpXWS6c6x/AfjHcP1YahvvF6zVu
oukxiFF4U7Zsm08LxTIUTgVAEg6SFBQ8NYSaANR/DTWyYz3bUCf+HeZKP/1iRWBt1yBI4x59SQcY
TNbX2xN1Re6iXr2iDD67TtNpEM0RTf+V5V8thJv5PqcvtVJP3c88hYgN7TfqqqELjEcYxfeV5X8O
7M+yC/UbPGmGM2ExZgVo1E2xRuV105DKZ9r/P02r+DPD0bcPQJCNJNf1gQPs5d/ECwgb0Y2tg7K7
3pOz+9ANNaaMe92homY8x6HhFAXcxW5rEl7qNuzDWAjLEsoeh74nYO2nQelgThTPPgZsTYGQHQ2J
udbuiQxkVBTZ+DxpDGw1fpp+XOfoUDPmUt/6IH/zAzyVw3BgPmQdjUw2UK32lg27o1oNqfyDgF34
E94RR8PKaaXNX5G0RBQ4wXj47GHEt3gAtfPffrK6g2jdhcIbXBuJIkIUfbZKDiCL318LAidqp1vb
atT17sFIqF0FoH0F04T8Qp+MwkHvCU4WVxZcChuAQxI/AvGQTjbTcWH4/34i/UPQQ60kGWCnjRFC
BIIrKrSchZuqrItJL9/3K2Yrv23c3YJrouC98NbODI0809jqv0fHq0nyFkiEEMFsWSz8n6p5fKv9
OKmVauN2+bXy1X+accTXAVMnOZD7MFAdatzOsl7L1H+RnXZTi+9P6RSjMPz+N8SQ9B87nIY65IFK
1EpOfC/RmSdqNtVlARFNebNnpsOA0PjPirZkiNLikYv4Zreuhr57Td/6Pp9WWRMy+rR0bzN0senX
pcdHn8YKUyknmXj/qq5G0FGjJ26aaTz8xiu4oT6AMP+z9EwMLEWCwvQjiNWp2Xjuc351aCH9tIEP
//xVYhAyaapcfMcLva45F+f7rv4ObHJSUG8lLluXSU5+E0J7LsdYSrdcqfIO2VwfUNKPhLZWiNyW
vgLxo0ghWf3rf2G9T+ySWVD99/YJdbFEMvj0Lakd5zRS5JebZeMsXzFYXGce7q4tFv+plONn79YK
9ApXL7Kl1sDhMO48peX8TnBCjcwk4ZOEmNvo9ZuYiqCPGtUyNxUHUrTgYLnfMGaN8B7zquRHBrUP
fs4RCGPREdjkH6IfpmeICVTvhhwD7dNcQUaID2rkTStiZNazATut6aykeMhbMRIT5qJ3rRk1FZPO
67v9bbWwu4NX7X9/bpGQWDjAPiChqsvVuISikYCIg03vPdyA/3qa0t3L854Fs7YUG7fFsjcm88w6
s/t2d0o7hIkSFjFmhIw3/lwtAqMeV1oxodF0D09Cu5USbT7To8hpwlah7wpXaVxeshPiTg7/KYg3
1ptIhEX5uWP2se0TDEx7bNukjbKzAJYFqg0Xx3hRwFH/SRXQmLHBGHgMvkLeE4roPysNEb1k4u8k
8DLvVz4GZ8pv3naM5KU9QCNZQ/FJMSkV2Ffbw4lahqX6CARhVKFtYEJclczksSdcQ5qVohMgfchf
5Jv8KaheY3ulnAQoUxswaTk07RCU9JwSrrO/VVC/2Oa58vN8yB0z62hg1+5qef0e1IeA6qIPCXtE
qN4++krsGtw/GU3lw1NDvNoivcZlgJbv/Jw05BBAmG5+QBMQy27CMGZFOXxsOxkPHvfQlTppHqUp
YSGRZPvK2aV6iKQrvlnfKH+dtzggmfee4h9Qc8vmGeGN/jHfC+5PApEnCiJh8MGSf4qKsWYUZFSn
7AxeRHO+0O7hhsK8x/nCOU5MFs6GONcNBSCM4TwWUM+wfjqdt2WdOUAIPYuHhCYAtL9x6y6RoCd4
lzp6hlgbZLvP+JwxlcC0GNhRAFWIgpf2Vuff08/fssNljw2Q4cEDCducgKshGKXqWTdFGx+OEs4A
BZ0svbLnEoVC09CgV1tLJDFAwVROYDiWDib2szz6e3Ott0IxqLzfzl1rfFLFSEb4gu6NYA3laIhr
lxZjWnSO9RRyKs4Btnr3G21AJUcP678nRYI3pjs3FmiBZp5p0gcaY+kQF1NNnWdj+4eBhLZDbhSy
Nh61yxlS00XWGVQQP7wlDd6SFLNlXjPohDqLGVo+4urmv1ARFlK3AF+2kEmHiJCEO0uaoGmj6pYy
fliYNJHhMi2rzT+O7i0VI7h8dkYL4sSRJ2pDnyzoaoI2GQ1fmiJXbX4pFS4g3hkBHWtCT2HnTXKT
u9GxhDl7ZxrMct2UkrMEoIjRvkQfhxIfOsj8LvMGIy8HvTtjfUudvkd5cQpGc6DgGkIDUqPJSoJb
UGqByKQ7Yt1Yw4vqCa5A46gFQxhq23m2qDpvzli/20p0JW2hdfQI414YDEP0F9kjZTdJPJVBocWm
xZ8SJ+vdMMnSP191b4N29ciZ36sBbo4tllehGmdsB0qFDst1rjH9AWhXKuc2NK2Q2aiLE4QbjjYC
w+RIlpxJLw0c3+0s3axGCFQ/kXZZDsGf1FEAVQEeTDMzkm0A6n1k/Qu8e1bZxrAe/ve3uAFVPh8b
oVX88mOoZC95lyrJ/x+XJ26sZOcE3zI+s2nv2a0CBMXGka2zOr0YApJEkGMnAE2lqbE0zRXcyF7h
1E9b7cZ5G29w2ru4keutIjpkLDeent7+SS+IZVFOyjVeMq2um9m2y/chXCBx8/g5dFMCtqeo8Tqi
r28C4YKkgej/ei9QQBv5J3fEAm/9TsERpWKiQ5fZwpAoLCVqmwegklIF/X6qf7F7Ky6HEoE7AiPi
TzdNobJiMqRFiqjHeWRgxbZ7NE2WcOaLcb5yMckN7XvWRH/+uOg6jr/p235oFmneidRPELAjrlYG
AH1ASKG78Et0Z9KMtFnRWmw0VxJBNyB/XNK/PAdBFALykHIyFutEZ35mLf5BcdxiVY24krqOEPCe
1YlHN/A3zNKEjtKP5R+FpbYBpQS5b7f3aMQq6LlZXEfilQTXsnK7QwAHevL03m3u7H1ZSrfdOAO+
cs4K+u6Up2Jqd6vLNnN9wsTzdsmqYcblX3dDe6/OKt1UqAMTeNmCdEwLkpHP45d93SWw/LQcZt7w
xcwhSv9e1e88NMnIiHjmAIC5u3E4jM1wPisRu1oNwuGi18RuQd5J8/+3bFRs6FTJ5zlOE175X5Uv
p8PzVW5EWaCcptmik+B3sycA/fp5Xq68jw3k94LlV3M39vkUOYYiJ8rGkLpv8KvWb5W4FAGTfgk3
XVSymrjFZuze+lfQJ/z2kZ6xEAuQtWXAz1gDWXHUcKtrpteCArkblMr/SLrMRE0vU/GWWJl5Un+c
sOEF3zg+itrhdRSKSPqrFor0IWhlJLhgN9VB/Yru7yYevd8R/BCVz6y8uVtL5JkQJtp9cD75mihF
EPyL5BogRzaGt70iMWxyjkkl3cB9ZbQBWy736klgyXbsgfnmKhYoWRbiONu7mTh8M4olKSzT1qP1
G8XUQSf7iA6kfXnV+pPF7IjMa6m6Ai08L8wqDGnUXkEqaGyZe7cB7GqyFRjJIMqkZxvxLM7AccEQ
O01vtRLU4fd403ptubi+obYiLVeJxxsSgtOaD49qxtj5LkYLPXtZ1SBq4OH8Lu7MDs8vhBgF/Xv/
auDNjh9Mzqr4Xvj93vBsNELi0fV1icUeixVEcmjmJpmKORhccgUjqf2232NPUyNgRwwuGLWZalxi
142OPcU+0xmKlmPd6JnUFPS5AppoeUJS7l7nT4PNextDls/zjNPFNtwk+UZXTpU3rJXjIWCVVMtK
cSfDBBBImtAnNAzQrItFCN1PU7iaxFEiajxDym6ap/FedN6KbwfI/MHqty6t8hIFVDUSg0t36VDE
cWN7mu5IT6Raj3BJDg47pmOVOog88v8AKikLqrDbT0GlIdBv1rbYaer3uyuvahRSbNu7FRwaCMOF
ye8EPSfmgh/u1MnRwP175Gxhu9qAd4A7E2p9Uy5tgQw0R6Q7BSFQbM5gD0nA03ZoX6YNJ5YWBCY4
j2VByLY9kYZ/gILh3X79hlz+5fhT5gu43Aw5PtjaY6H0kpclEIW1VJ4z6Ifu/+gfgvAac5oqWvZU
hdLe+y6CHJLg7/2JDiOlehqOMqbOn/1Ge/OJAKl3HjbZOE2k9XCe4/OBBtHo0GNRCc7WM8n81VRp
eApEe/ZbP/UhfASDLZIEnOb0z2ulXINU1vgLFrtybPocPx3v2lHBJKeKbyv4OMhofcLGEK6rbjjq
5bKNFNSOMONLvf8/MpQ+2m3nqTAQEdj7i/AOyNU0cKz4iyzSqon5DUh0++LmbJS7opD9cnQ40GbW
albVJnbqmRmtv3KzO6NtRGj+zpJJ91RjEYgcUOPSmH/gSJH07IVsZ+d9suT+eEnDhDwOXyVQBVH4
XB2VdumvvSJNDKB7FkOrEZthJhh81agBXgpuvsi9TjzvtEat11mBpeE5rwF8yqMlWX2KLXM8jW9F
gZpZ1veJtDU1SvtfICAT/UaX1Wehid2qpp9HVHzu7eqPWXK/HOOvEG/L7jZfJeK40WxS+6WB/bXg
Pikz/qzwPG4Bc/IfATLge5bCPKCalyG62qR7ibuz9rWhqO6z759RLihsS1N4g850fctAOPM/7z4D
xWL1Lyh1Xx/5Wk3o8AE+1yDI3zECcxgVhG/QqxNMD3wvC6m6Mp1ReurJtxozCteeroeBzhU0eLsR
Z4PqB2TX33bw0xn7uM2diI0VSQLDUT08BgQ4cwQ4yRBIv7Sv6cSyOQVJTaOeb7r/PRIGSLiOfYVc
Z61eebjply5UW1P25C2F/wWsZezBW2XVzD/pbzm0FEafBbCVWk7pgPvnA9RJuPCtWVguiiJ2gTFO
seqCf4Z9LxeXCMS/duh6w9R+WjYkbT1SLbQN0Y7ID742NGb62EOz1Zuwzc9cO0RgHfw8yi8nwmrC
lzbImpeu1vXk3lvJuQxvSy0Q8GMqAoEtHHF84hphnVO+FhY3IrMQaGyZGfUURpovIa6Nb2kiZnXi
CsmKfj2fRklMSKU4fyOJlRq00RDS2Vzqj5zRJ8Nuqc9z1QWyzr9W3bBisKn+m9vMMuv9n4uRxaEP
05I5w2qsA9CG3wwMNroRUOfZr1ubug607iigZVshfhh3Gl28F0MOr9QBfCDtKhbiUsFgsoTeolQ7
ce0yEqWc+3uA96owhtvLUA/RGbY/tJU+pPeWHW9b9O3SY5qvg4bN+Z1TbqjTZMY0geaV66RfDrdJ
OaeX6qi4dASSF8Zk+xdZKbg6eGGSILolWRd9b325jD8iouo4NTEzTouEsOGOpJf5eqXetHHKXWzc
H+cwwGteiCtlZSueX5mJUbnSdJIBH5CFMXD1CEuY0kI25IkriRXUvyEB1DruuKoObKKHOTTf0F8T
Qk4rhQxAQoGQlmmAg5NpvDpEiPZiHKdtbhHFQ/JuWrU8Mlvv2CTv4xpw7V9+qGxplo0evo2dSCFn
9rdGxsa1853S3ov2LYTvs6CIsqfpLahdBDjZYzWlPQkrGUWLo+i1BIAo6jC3PgqxQ7j5GK8xguyy
aPQ0kl+PT6CSYhpQpyGhjQWV0JUy3taktJp03AyL82+1CeIYIOJPznbqNVila0TevE1/tgCHsMP3
0qz9XEVR8ml1bTzTqz9frpEXWeryMdMAV5qCZFcYr5E23d7aPiZ/4lw9+xbp2odk5J3V6B5W2njE
cAPiota8ibQs+bLUigs/WzUyxAVqeuCuMAIU1jqqZRDjOUGbopxk/06tzU4Y6u5aTQ6Eq5sFstrD
eXG+vORXxyW7Oq2w8iwIVD0l5ygoZB6DA4i/ZwZxOX0Z+iplxLHMjKiXJ3jPKDZwcEjuYGNf8Bxl
kc7GLyomvva9ENtOhhDI6A49mU+qswRt1hSb/rXNCjEXMzPx+MrZIxnY6Cxl47BZC9O0vWU2VvXR
NEavTRmbw4/SizSrFqshY9vPxVnViZGuWgtctVA9GgHWoAWPdeOIQA5bNgz4QIKm/AsqMgjVeyJe
aM8y0xEV6aNp1AZi2QOeFKhr1uYChxG9aQEZ0FXDYZ2MuV1IHy+LSGyNQio9nDzYBFnZ8u567qis
NUPw24bpQxQyVwLfRn4mFctGWpZX/bmrBfsdckBX1VgrRXyyH3EBS9iGCuJ5nr3ic2Ajn0eeloLs
CI7Fg2LVkdx2z+d0fo00v98G4QoeW75etbWHQDJ7Lhsmgfej5cetNSzBrtiiTvWi6tAE2oScE1Os
VQsI4tBoJQS5ZrDX3RuMA/u0nx3A3YFM/MgMqIpcp+21eWBLAv4bGx/35eeuaSKMRbtSAr0zJrrj
sH0392HR+e8PXXoLnNCO2t/wl+yQalevkNJDUkBfScjDNjS9CHpyTij50tnXYf0c9jwyC1//QLnt
nrZYu9lEdUYySyO7fof/QG+g7hh+JFMevz18MDEURWEeq83+f2U/f4KJWst+A+td7lhDj9Q2OKbx
2bHb/VgVaz9IardblA4xB8ZmGI+DBaU/pJvXBEk4HOP7/JazfzlFcyS5mjlGwKcAT2ylXK54nggu
SXhESKhvbs2dHhkWmw9pSTSWE6+8lNj1eV4XUmX829yssKR5nRMQ7IjunVBgTF2F1wZW5biP1pBx
NB9xYciJljL9ZGrtbQOrMO3YJN4xCuuBgK9S+VOyLXfaBqcb2qXHruNw2PXZqn36aJnYSUaCYN9N
pKXzjzYWV1KsWwxaU5WaGScCIlTvcjHnInYL+VrZ29U9h73cZUogY4m/c8KU/0naAke7P5jwJigi
n6eIkkoaFSWKLUViv8jjfUD6ISC/YeMt5G/VPrd8t2HJHCHK8sYWjOrT0/rsF7xHkiQEIIAFiF1z
3KR5ji2WAx8oGJaSGqXR+dYkcol3Z0tGBeu9ZnjRP+Erm5or7FrL/if8y9nP//Cdff+rZQonXZhQ
cCQJ8QbF7gXkk6SpnLCZ35nxytuWDzd2wmwAn4vc+ZoCJFB097ugssrr3/yfY72cScpK6Kiv/pff
znEoj9h25O7ipcN9GWT0n+Mli6a/AdwUJ+UJ5A6G5oI7w3FFMEjkX99ZxmLnHG8y9E2+Qvfjg55h
9+xx55qW5UkFpXuMYWe4YnQtlrs6rJulKwjHGiJOabR9/KdqoB3593AQnX657nFrSXNXQXW/aJpD
XOF6FHvwZZ0IOpJCZEivIYwkL9mqBR3V/7DDKLmv5wVw6CMg25oNr3dslGVBdceBz9SzkrOmN7Rj
7vMd1JFEbTswkJ9dlrDKL0XaWUue84IRdHU95ABMXYlQiSxn65oRL0lw/Ft9+qIzTa614r2c7yRD
8cAd8MfiGIMB7oB6a8hK1nB8aOLXu2lGn0xBIVLB7D3iNjQFRy5UE1/jCPDpGm7BceDBnAY6TAYB
w6/Y6Byf3jSCC7nsPh0sWqIFk0tBSyZshRdQQiZGT3fF/5sVWAAKredyMtIjPDHMoQEDqwou0U6K
nrSzWHFCmgBq3TiKQ3nVCERbBvYvjKto9PZOhLpSgOJbIvweMVnsmbr77O6BnFp+ILy6Ke5guXtS
7G6prJb2bYnlIZnFuuWxH8efjOKZASBaEJsa2LnSETJ7WJkGgnVAVrz2hwOLaFhRLdJA45ZLf9Cg
4h/AYTycgpkz/vpT2SVWsyJe0JrvJbOTGn+VDsarGIoW2D3Y9uOeYpIqZeGA1NqqKWZmc1W1JDtW
huOufGmQJmki+Tv0FYLP007bl+AbiJ0LKhPi+IUAATuK2JAjmY6VPlX8y9YhMuqxC5BAEzxc507M
6TeQX/zgnIifRv3Mnl91kW8pu6NBQ93/nFINb5jlYjydZbxlybwLIDMgmhSiqoaGRGCse+7GlnH5
fTcgAsVb0BBYaZ2JoatTsPbeLk0t9Rv0dnIl45SHAZABErmkRfVSU4+9XdFxMVVTwWGxvuQxfffp
s2pb3dqjetmpuSRnTPZJlftjZD5I4rIt2gdMlxzzBQX9d0zn3v+wP664CnDfloFWgUBMSrPq6jhp
+7xm8AMAd79SlJWMLWhZG/3R510FLIjeo80KEyMkfXbaYOtxtkexGugAlnw+Bt/bKzu0r5awUslb
uAxBTps1OTwGnRkgZ25t7CS/GjNNy8yAzL9wSMq7vNFB4THtwCDo+c2H0IMBZyM6P1G8zcITKNX1
ZcpJkp3W2p0mN4a31gamkr/XLeqTWxicHWdltRQSwLL/UZzMXL78Uito5ABCwv2r4JZqy4uyjDlR
UdeYOaq+z9W304eHOSPD7t6mIMFTAT9LGPSaoSILZ+L6J8s+yIBHiSQdNNscN3MqN4Z1QsEyGfav
ZPzue6tG8C/3sLiH0c9IBQgrh02AAfXMPC1HdPJrCz2fN/CEXAPeTxYCzgGu1/2bgEqnQuC8jpP7
t8MPS2HFtWIw5Xoh5NpyXbbUmLss7i9gEELqkGEnXvcjDD0HdN8ZxvBy4p+zknRqGfNI5FglWs8g
h2W9kbKBGk16lrTnfTT/NMho9Mst19e9BO8Hq/v4g+g/DXxwJMCJuDsVqndd0gP17McX7g+cCXdM
YBAuAwKsmpWBSMpL+/3bqm8GJPjwNMNhWbqIF1Vgyo9vaqdxjfuxFq0+LdqY/OQbXoQoWHjW92WM
posaFFPt6VZqjsBgK6bbKCwTRtY4Dp/L8Pm4eYkER6BAd7t+4z/nBlfGolXp0zDG4ScDiu2Hs8NO
hu5uxZ1bYxnVOkWzqTMnxg6yJYGf/XYCbMORrOg5ddCUsDyUl46YIqPNjLL+fZpALblQzylgT1Fj
Yy8CkmpazBgn5zjf23QcVJ7QG8AOGsANiwAvnTyYnzOs959ky7DMvtpGcEMWzv7E6EJUk6SI+7Wu
z9+hSZo7Jz7AuF1sQfnZY0eSSGtqb9p5RQ+1c1oTnIavIkFKftRyBWHhxmuQFfdDQ6QFX925iFEu
LKL/rJH1NgY96/LR8eLwTf4Otqloi9Na07HRFzaHLhDH/LuQakWmbYlpH+QNrWxh5qC38csb8Em1
mC4O7ixg1yoRWTC9VS7eTYPIt/qO+n6k+M1kOq98972aWpzXNftoueuImU6HdDfCoQh8y7c7pWn4
x+JcZuqOrOnZgbtVqxQgOseL+c8xmdLj0moRDWkYxgGEvkughIhBsMvFjcEw3FAEG6Rtv0Z1c/dW
T/Zb3TSfEIMbAZ9p1ZgUZnU95R3mR8g/f8gcg8yGoTReeijtxaAZoRCz6OskpcDZgzor5P9G2zO0
IiujHYG9qlRdBG/K1X821L+yta42LsSfoOSuNBKamRstwaIJ7V/tUCVD6Ni2huiHgvXJO3RSWIxx
00oZttTc4dTgGsl4XHvUmZPyGpAXe81Ip05IheDL/Qk+TBGSmbhNxVzA9qTSX6uVabxFL8LZz/5/
MQ2rtWTCRrMSJ09RPzzlPgFnEyW/PPa2HVsyc0e5WXyawHyRO+jzcgEJK+tNCpOfzmx/mYW6sQAP
guBXr0O6ikZUe1V4Nnb0pLP+MC0TgdFDQP4SChFaKcVSZRagDrfiqfK8HcGyunhpx0pRwheS96+8
cilQo8X3EkNBKbTTL51TxipgAV5jfUi7QHdiunOgu9By1qiqS/d2Y5lqTD6nYCIdTTLbm6WtHzrc
IOyvRArNg8+M+4sNQubWUiPYcH53DOYfhm3hJitWfXOs+CnJVJbRphMhNq5BfphqrIjRD6Ia+Q09
ebiWl8yEgXGwHC/8u0WMroEh0UeLEqguUCUyYvpWkCtKVns9ZoTMZHJYwIJGm/XE50hZXspljiWt
qsqzdnHPOYfgM5zp0HBEzj/xIlFmPtominarQjFHaMxrECvYzdrOobSQwD650xtoB8NCOcvyOQpn
ZduNSb6LMh1P6R45tNgM7tc4BGw2ojSSPcAILALGncT+mrnBZ5A96ZfMPEVWmkr7eLaYlo+bikmm
z1o/whYE7q7rUVd+v3gv8Vc3z71+pTYT6UmE87aih+4FFKeApBiuEM8VEp0p6hkN2qJkilGy6FoG
L0ujTinx6scxTA8m0GB9QkshmGRk+PeWneEDTm3tZSArqomXSwPdOJaJujabD1swCDdnId6T2kci
i8067PP2XBjbeInw6Jbr74VB0THoV3PzIOp4IpFj6/DnoHV/ZiiV2FaMSQGLB9GU909RV0EZLp6p
WGml6YG1MSvjnouVETrbC0j0EH872uY7kND92+EfBRQ1ecfZ0G+47xNYMJlo7LddpcKtQg03xP9p
dUJWPncGuMLGrP9sQbI7QkSxdQSOVsOeoJEXm7SKMRq7UtGeW+nylRQ5yNN/tyTRSl36TgDxaaF6
M0Qc5KMYSK1prwMeSqy85SlYhBXKA9BOe3sGJQyzCdalf1+1ypu/oZsPqZ7jLkKJ2BriRMqdrLzo
U75/tZKrPkr3ez4o+/fHZxabprJ0hSz3ThSwjt+AGdOyi1c8OcJHazcMHz77ETMTx6fMK4Uj92kg
JAQOJqy/nsRKVqFhSJmC7uETP6HLCRdmpoZz6PgDT3lXL/afO01pOoQ4aPzYb53JGnRrMSLa+mqj
T6WtsRUSQwYpDUfxZgfzVNT/stQs46WEfgPjzZASiXOcTGjRyY5XhzI2M4NDvTXrzCkrs4K2+gxv
JJKIIY+tnMPTlw2EqqHCcsXWVHTqKkwRtqVOLe5H2XmMLhiI2LTrY7TfvFclQc+dfYvQIgGJb8dh
zdRJa5eil8VLX1fTZd3JTom04wUvQvSskhWUDa10EyYEjTIi97gVkD9Okni+e7pvdlnh6v4p/PZa
GjRi9TCoYYVI9QjxNzC/EeBDCIOcNLVGY82jV5kkmaXYe1fCbAmc079pYNIeND1g7+jPLS/M9PmE
vCeTPX90qLcu+f53+GtqvFuemCjeNfAWZQAmsCflTvrhU8uJ8ruwRCm5d9izy9d0EPtZ1Zd/SEYp
cDQJ8V9A8Vk3n+epLLymN+NiRP3Y9plLrqKUZCT0+Azgf2axt+KP67m2GWQwmlG+cfAMLq73wf+y
fSZxUkd7mn795DiEhmAy5hUpTfrJoYuV52Lny+tAfxzRynCXhxEjrjJHJ20DhZhye0t0nRxF13h3
eeLZmFeUjkq0Wlop7JFiiqYatass/7FK45nbZ1uYHA2oaP9Rc0Ig9sJVhZQVXdQjBoZkXjhbF5XP
d7gLFh8r/72H/qG0SSVyUpsep10dgDUd4Bc1/MIV0B7VyFGoLo6bJovGVjEdBT6Im/NdgC/4QCAY
mvz+c7+Lb9xKyizcFg9ObQjguy2x2i4/NjgDlDqlUWl6UqNKsnlAhasami4RCZOqgxm+wVLR7o5z
qoade57u/4qt4HN3PRjs5NW5yHlFY4rPcc0irxXGZp0cHnZVhXhPpYe+ieXLxMHesgkChrWtfm34
pKGafbC6Nu3lh++EMVCjnfdAnxAo6VQK3vH41+dihhSKORbThScy9xVUliLKI9B9U3Ow8TYayoPg
DTmTpYvad+TIdYAwn/Kq3XZY6T04RJ3R5Opebnp9xb50EA5dNRVF6Rnk2nVkDnZpVUi6B/pr/1rT
H6fRLNdBczM/waTyC13fEs/tNsItAOFtXA5AQNZ5x+m1Kehx3efBPVbumzwFT4n8Jh622kb2sH3h
B/NEMcL7+MTr8ztnwtTFmzEpPEjIhb1TcxFyjo3mzMBSawj9UK+lDf0QIc/qk7ADvfxM/I3Zlr/H
M9nKq7HPGBcYxs3jtoWkUH89aawl2dAZzAxz7YGbvCJm77jtPZR5AifEGACtAa88SP2WdjiJ959/
u4u52OYeEEjYgWVEnBwB2dMxyCWPPU6OFCjSHS2mRZeufmFMnocJn5bejcS0dRudbr8CAewigP7O
ZQbOiu7JySM9yGHNI2wY9B6dqHOXE9sMV2D7Q5kfzg+Gas7fxc4zl2YQTfgYV7NxmQ/QK4pftA0N
iHMUz4PKncmBE7WCeuAnx+dcW/3hrd0ZqqPSm4aQ0hFXlD6VPHcismedRMdShAd6LYICGanpOuV6
zHZgNyDsbUEIg+uBhJPgrcP2zaB+vp+fZQ8zEtzwZEr+vgchLBE69ivnLO/MV8AnpIBWIced+Q+C
nvGMqDoW+fQ1V/3UCFzyuYeCXNlKE0Z7C+0BQ1podQnrymWtH0n4B+KHQJ4z8OKytwsyX/jIFHFi
SVbvAe5DE60D+nk42ZWaBVr0C48e4o5+QyvTcENF6G18OR+hSxdimJ83irMirQLindImuY3znn38
pOy9IgntaMERFHorg4V80vxsBOYAbH2uW3RyN3B+XhJhQfx8xdg4fW3HedhSTD4DnIbyEPLG4NaI
xqVdgNu74iVoDUA90jVJfllrIs8XjnfpJTsvLH82hmaJR1JP7wVNIuH9sXZ1JhuVIrbrnDgA0DD4
RmwlHybzBLRkFDXwpxYLSWTU1dyms5m6PTuTi5LvhZDa+FExM7RRTMOFfH7534isENUTY2oOM9VJ
w5b58iaup5+TpgLT2k8e2gG5v+ApDxQCCnWpd7Fqig7toGZJsWCqj03yo4GayJS3ibfwKYNzE7jG
3fgVqUJiE71qanWnKXk6I8YkrwMfzs6zvEPgCuJhBRDHc/jefquH2A32j32QRzAfZKdXsP6VUtMX
OzoCZA9tTNvurQXFJD4WYVGs8Xu+rNTFIh6QiskSdbzxFG3NTmKTBSGoHbPR9oKaDafzMzjE7lYC
bKJAWmbZg4Ek5f4c2cOXNfg8tbbhv4Z0q0316e/0i7ijRGinpKTHTKRa+Q31QlOAfMwn5Ur6uKrr
Qi3oC31cNyBvPEPbM4hUyF/SbpJ68frvqoSIWgeYP3VM14/rmkSsSgNdl9erBWm0+5WK334dlntX
xGtRIWbbekFsFcXwe4tu+BDat0cJ2dfkt7V3bEaGax0gTHE/drezG+4m2DxzVC+LkiOKTM39lzSc
FVLRgs8oQyPdAe3Cu0rjLRSYrFDpr1jJB9gyhriWn4mwHCKlcrJRMtoluvZLtWyaN7Oay8JhH09e
9FlLFx8Ogu90w2NG6EK1cDj6RtuunnzGNrTsXurRKF4xmVpGbUxkF4riIDpY1Ki/YIAjBVNr+xQf
xFBkZHqtYlB23q5QkSnfcwG0+NoW9zX7PX8Bo5UHMwn9EPjsvHQ40TdBnSBNXo1HVaA6Hpfd1weB
pRHmlpMCbf+cIgTZ3p98om28tMfAbkQqZ8iHQphtwpLjysIVI4Uk0w7G4uJA1gEX/KnXrSkrpJkI
VO6WgfLqa/qBxq1aJS1mOpplny14jUSJYk8pvj342PyijhknPM4EZOiYTx4M33h9w8NIfafXooNp
vdCsGiZi92WemEQuH2U6g5UszxBb7jCWtw1n10Rca06X2AIaWgXy72ouJPsS2+sfzqXSSV969wgP
+rvp2scmsPBdhJylGTaOTGkXLLEjk/z0KHbUmkn+TaptdPGFm01QZW7zaL0HSf3C3qvjkaPpP3G4
jyP3zFVkrjGTbWUNyL8VjxsxXOJfWNA3tMQjZK1a1y7cciJVXuaqpFvp+21ZA9Tn621IwKH17gOo
LEtnHM2lJZemEILHgtq9Pawau8+/ryZxaqdvQNhzPWiSkVY9mTfrCBvFGoINd9TDMdIgDQzbRe2d
b1PD+hcJIV/9gZ4n2idjiKh8Ds1KHPHV8fMzHhle5pQihHCwAARmDwzN6dTfEkMYwsDOWRNa9E5E
1YhxbjXS2GZlJ/CvhIIgQeXXR743duJ51pj/bM9bVHwZtTlczq5Ip/j2DZOwlBEmjl+gWqkqcw3G
rSNOZvT9pIpS8awn2aEytehiznS9p8qQGck43+kRyoYhU9lghyBalRkT8lN4CvGUtpK7OyWDkW/r
1symq+9pKe+mZm79oFCAMIv4pR4OcQMu+UhuQyB/ialSiP1KFKMXwMmSQ+TVshdEUwNjvQm3pgYJ
Yx06/7vRVHFpmm1CvGeiLes2fhEyqhKqBZv3BuluCfK9nxjGzvGO4h4hfc3pzRWuHfUFkxKYtXOf
0jRFJesMOTrFcPSOwARAnbN0Q0TpZ7WeiITtY123P7JkpC5oXAMHqboL/5+sw7nGEQSbePM1E5iq
IeuMmN1mDhbRHeDqFCYEgMNtpjI4k3n1VT9n+cEmQHLX5yvSt11GKkSX7rujARN5Iob/r2zVjjX4
1rg77Wxzey7RLc9RYA3PJIT9TcC3f3/CNkcrx8AwXeGwRdAZdjWNZ9AK081zM3zmEnK5JpLhfuq+
fn3WN4Cbwu7i6AZaeODX2k+WnOf5Zq1MFZMPZ+/JV0caPX78ktnSzYpToYNc7GWnIp004blFiNJm
HwzvfKzeydYpj0qRNQBqDOSYMwlJO1jkRsgqaWPCKUDgLXsMVAbwzD6KaXozrpjP4ZFKW8W0vr5R
m91em6Uj+lGELVRrzByrEYw31jBTAho5vl2RcFvlRnS9axf0aImoj2sSdUGZcTF7lSBDA0MX6ZdY
gUQDysYYtsr/oXy7LIXXYkJVqpI+km/AlUiAl4/G5x1rFvNwfQjf7BygdAVIq295zce9qWP/1zjz
/g+QOJzu14Dd2eUELcZCLhL+gUsMLRmPiimFR56OkSrHg1qdziUv4aJ8bSTjiwRBd68qEDfgfVEk
GeQvkDinUW/CLmSQSIUd8d2QFtQK23Xa//RV0Ex8cXSx8CSly3PbGrFEqhYLTYgVTALwMDBrFhke
YqGqjkNjYqe0ZMDdxRtQ1FMq18IQOYBd55rozSZi3ke6x11Seot/7hHRkgiqAkbzWlZ6b20s9Njm
3gJRRihVWIYdkS+o4KmvQNg8zHM+Wkvq3UnSXyxEy8GXBouqEmqCfxogS7keO2V3EJzWVXApmRms
K0wWmAqOjXasj4XUhwzTLHQ2m5PP5DY5aq6qbqkD6fhO42V06ZIXqkAypX0QhEXRv5s/dLQ9Nexy
f+1E3059AnZfc7R2Eg0CkCP6fnj9FUXPF687myW34H+VelDfKguf223iR05WezZJ036ctUrWR7cg
wkfRFEWqB77dF4gHgFSSjAuI5tPnOiUyzy8mKnkwwRnIk2FcqvF75kNtAeBD9Zimuc5z/4mOifgI
b2i4/cc9sardyY4u/rKX5VMOde3/uHvG6nXtnUi2e5OeP9Subi2CAd1twt79OkXWzQscQ+9V+Q/M
9mFBzuu6l1Lb8W63e+WVOXD0kGHrlh8BoJH1H9FqHhSn91QswFrYcABtFvMy7Eb6pf6Gsp6vV3dK
vSxf+15UiQSxUJs3SUjmTWeB7Uz+jccHVK1ycI6Ube3DSecjFRb55MHYES1157ZC4G3Vrp+2r7/l
hCJuHp5fwNc+ueLIi1N//irzc/dt3gjnBn1xbJvxZjvuxckT4vY8V9wMoAPvPx2nsGGuPtyGDAVh
Xet2s4LIE8orUOG34JGKI2p9+d+MYGq13sB5Zek6ydWZoS/lO/06q1Hl/cLc08ZwyqtqW1QUanQb
Xegxx2N0zuI7hfLLnRqU+QmW6r/D16AbGioQvnIxr3A3clIz5bTetwMU/6jqkb/1KXXQZqIDsvSM
0WvcAijbPWcGLOF/0ZlcUc6vEQjhxE6h2it6rc98GaKs/QQ+fnDk56m8kRTaWMpStDelXnDpvkOO
M+v5E0aMV4Sz/AMwTmFwPYIQ2aY5Nl35e7ILk3bhSnFAxFPYF89GstlSyo9NbkW5zDXMXWE6EVBX
nWcExu7HH3Blaj9XIEEjXlBH6s69zDVsVXdZ2aBXZbPl/MUttV2JpBh+rQdRZe/iwiXvXOclcO+9
9Tu9hfxgk3Pyeb/3zxHq0+Z7HXz5wqcMLn3ea9vEeocYGLBb7Uc90rW5RuYgvJ5SbkQtybbL4oao
17XlZMh0mAIMui4LBdqy1S7YmBt/2zM8FcsAppcbKUbEx2yHMxVgygzljJvhGMxU2oZkaLwDKMe7
bwaPsLsk15ECY1j3mZ5U+XF8UZicYznp20QIVGQqufIq0yOSKDlehVTbFRFRFt91uk2L886ppmQl
5WihQJ0cg9a2DLfIvdg95PPpuHN2NZWB0z8vAF+rEm4qgR6BpzvK3VNUzVpsLqzUriaTWz38sVsh
uuZfavxi6r+5xlS5l16KUZMsqlBNlIB/FwPatleyQsm/JZ8xg9xekrffQfmHIUaop70jJbKE1t1x
0j0Eyvu6Lc3MBk5+3yQujxPOffg89W/+jLTUT+ylUpYwyYnDzm3HEjOcFvxuS337DzqD7RA+U/dM
54gF8KZwlKhAFkj+H0ZV90UMdpF/RN6GpAPICrEbeZHmSkf5nZxoNJh1aeX3oLhx9FzP2DXtYfv/
5HgSQdaPKkUQb2wXuud1KEOeWuDtUNZODoxhFypNayuuRaPXflxCMr/MviFW2Kp51gI9XFDcro6A
JarngPqCzkrSotiLg0Kr6k17qV0FbK+UfLxFanyuGObeP0KP2Xv7Aa/3xyHG+Y4Qux5DE2dTGy7C
61IhkaKIc+QFOEgbqoRXPud6II8cfnToU90Un4aA38UaLY/P5j+DfmbCppZD26Uqka+h5vIuiruL
yemFAhkxiUCyPCVzgwl6rPv0p7YsWQeBLLiN3L8A9YcpgLYOdMubZl+kInJ3FTHxQzzXhBHjMsLu
ZBgUGMu5fuk9ERAGqwyNFfaFjz/bCNb/+jaLD7YTwS9r0lbtiPvHzHGXSpGo1fctpSSo1Uli9FIo
p35DEkl75lmc7+k1h74JZKlFqpCebMBqrSbZpjKqi1PObwNfjGP7+oyJqhYaeyoM009ocpZRJ8hd
ba+7P8TFdSZxE6tbWchooFudONQN98C4vZShTLwhIigA5SsEo9oFS+P3MecsYK7nwV8qEVjRq2Fe
b+fH0EPo776LrxFk+LqhYsPNeth/FLBXRHLGkxMki65ydalqR8ogacBHMhcnxgGjEJ3Pf8J4tQb/
rsAAJwj5tBCelfp0S2yxWychlL9kvy9I5H3l8sy7vfrm3ufVONvYkk4VBePUkb6ypyMXWutjIqZB
i6Cb+6TrT8inj0i2ro6CQ+pIxjV3zPseFc8u+OJX/AlnhL+Utz+d9oJXv3TdCljXIHsmss2SPM7q
4mbvNm//ZBX6i4JEVh4zDBwH9td/WPOzNm26KjaMfoxGR7zQWgH8zZCz+/JXFBbX26YOu5IeXe0G
SGLYNDBhU6KdTxTqDf+KnjAkK2wS+Rdk+4bFxdfZCTtgLxjf5ufLyvYmgqYjbdTfcC7M3dT3w3gV
dNuzsnRVz/Bb/t6oZ7gF6dT0ZIfOEVgeqfg8s9ys+wvBg/vkGN8IlNsLj4eqOFfQ7UNFX0x0l1Ug
8SbmQ/klzyv9VmXmqx1psIMIi3HCiHYNqRX73A4+l+Y76hl0Hxy+yJtBFX7Wp6T5IAo6oyU9OX+T
GDoGBx4CfiLH4+wFYS5zrOZPiaUEqJTezBzvzTJdbhEx2ySLLg8dGVbtKhAt7USfRHEfSZMTgVjf
Wi1wEef/AVTw+s4Ohpy6PyWeynxs3WBUr4gjcsvII2bEinT2oCyuu7ha8TEono60V+PRpMqxUN5q
P1SXDUFV9V0FB1lCCODVMNsX2Fx0kX5RuxS+b8dUEtoZYmiBBNACnaVvBES3v2Zr26eYxCa7mIal
Ly/JBZ4kzTI4Wrbx0JRulwjzJMFrZeu36bXV4Q7GIM/D+JEiNbAoE4zvANJcUPLsw/Ql3bBzywiW
QJ6+VG7Oe7CDfqcQAtvk6zLdL7w2YgsMmy0ZWKFSuVA//1yyfociHviQKZaqCUeC/uLs8bSbxvxO
b14Yfpv3X/PniQbuixf5LO+4QcZ+Yvni0/65YbJrdNxRKWYBsFplxBDA2WtMs6wf/PxDoKGsB1a7
bwFxlv0xegtxLCGgGX0O4C4PUDWogmBTznCt4C3kTuRyqZdt+th/CYSSz47a9NSjO9j20Uc9SGat
PRC0lFxt/DUpKPmKEK5PP34zshpC3ZYeYE77jpGF4HoE1TPecrWeSWl9VyYIqoXm6du7VBqSDd5d
r8y1t63HWBkMfU22nkTKjACR3f8NaPZsIlmzP4F+3b5fdXiXn99xepflcOmw9Flc63Yd/zK8ezOQ
T8CYXEqPCXMm8BInGSDXmtOy6shbxXaDYMqWdYupI0B5y74BT94Ia9gPU1MLAF9uDO9qjM2TI+3A
S9oWuvbDZ9ZagVA/xR3B9nLwz0A1IcyTAzYf6fQ4FuV1Q4otfwwwk0lOBXZHSDwyU8eEqPTJzUdk
IcwaBtt4sq5vQGyzyfsL+cHeZ8KKOlr8BtB4BT6XQKKmiEE5e+QuL5DpIZ9ttOJDr7u0Nap4hUcu
adHL9bmOF0rw1+U5hu6NPo/3bpaPNP7Nlpz3J43BjLX+swwwy8QdUZZv9afpAPH+c4Jwt/jlIJif
EkdLsS7axnHbEt2wHWgNAGonr2pqyks5uWOlv05+JB3IOyyrPuXr49GlgOM04dDXHo8Iq6wLYLiI
kF7hySXjTL4URTK6pGcMo+c/gBgcJqk3cowPI983bzsHxY71+8JnGALx7i8ZiLOobGsaXDVYID9U
o7ZpLxO51oC/WuQ6vLU+YScLeBU735PNJIXVBfQAUyacFgRGE/LWFphkjjn0jj67LqVQDXGz1VvZ
SZctPBUcBZSgTUbOhJRUqmv1rMjPwnsE/rPmy+QheTk79ICTQE2Z209W1hfKuQ51ApHufYNU7n9G
YQOSdP0w5ma/UiXv9f8lT9A9v9Y3Jl8BHOIGB4seILjumhK1Z7PD77A4+N71+B3//gBkQfD5nN1n
qQqfA04KGLjzIY+e8YiWUVzZxawpx1+ZU8/y9tt3IYGTw6wVaQYWJ2RwW9L1Y0oAP6QaJK8vtdKp
Iud+xp6ZKv1hq8Cn8lcYOzEeU/7IUiFSyNNnLZrPfivKtLq03xICL+H43Pj1FMK7ouwZlpxa5G4e
2QHtkzqgB2oIUL9cKaVzsVXps02was6idzzkxiy2n+47/Sq2hDLGnpTIBfFlTA+PAwJTB55Zs3/G
tavv3jLz6aGd7kEpxOzp3m3nIlYMmhTm/+ucb0HH601fj490uCvlJOLxmaryG+vrkFHW5i9TbxEx
U97oylsO1nwnFgnN0MuNtEnY/Dla67WLJ7V9E0t8V+XrkKx5Wc7Xvqeg8/wGzmrGrk73tumV+zA+
rqDQRM0eybwPXWHT/b9kcPrCdcODlTfSY44yH+hAa0VwiJjciCdFmgT87Qj68axCw+XN3gwtJOjF
tefg/chWBdxXzTLZita5le+fN/Yo8pzA/AsfxSspzzroE22+S0AQVoDuk0w1kuQLs+0Eg9of4HYK
ZFTCOnokYIuhNVZyLE1j8/zmpYXdHYFGGG2Ec7okZkhMtZbWA7UnKgm52/qlNbQADigF4UO/kBA0
1HDYx5/jF/DKvivNiEsNBRKj+F6ICHUuq+1yR0GLwfNPwDPW4VRrWGnHBvTzFmpWC0XFP0mdfhXU
HqLLI5V53TrbF1W3PgeQDRY5fMQN2wduTjPHIfT6Jvs2FLFB63XLxOYYt4U1aOoJ9phVnaVdhMT9
TWITYbLd6BMQkyyBgyGAojIx48bA0dhe/wmqMln4ybkwCHMPF6oo1CIviisC1ISIt+iiWZvxZ3tV
ep+nzXZOjYQR2jVGQ26lNCIDS0BJoGUxzebGPiacmdmE+sbQh6szMdnaQBeJkWk5C/kICrChb0Ey
VBGgjTfPGFKxl8UBH9GrwUPPqdwj/rUdZnDLfPX0J/osst2FjX51dPQ+GrVRIvn2iO8C1cZDlYDM
3N+BBMckGxrKlLlqRNs7hpLhQBMNnwoN2eRvNkSULmBgLJ4kFrvJjMIqdP5YYfMggo3hQX8V5zhW
/t4kZbNhxQRBBn1xS+ug0fRsNeUspp7aOysJsHxsHrRNaGK/c6SBtzQE/ASNi42Z82QCzVm3JISz
K3ogKBHLNMW3raEAm/VWhAGjaEbRVG2axqd6qEiLuXeokSdIzrZi1FqCI/6EVBuPVdNKc4Qbf2tp
tfT6FaZmKTemlZyaBQ+5zmPCtpRemfwS0OX3/G3xKN+kk45gTwowgFgjcru7XYighzjUQxBf5lGA
m8nkyCqPGQTQOVFVzrc5ZPVR5VHiNmwYHpbcQp+JbPZgbjnUM9s13M+38NH3bakQZhtt3mtkezsO
hgA5iJgbtVV2WXGGfiThOr86UtyKpwReitEsUq8ACToNsGRf8v7SfdUAR0uPHVE95K2fQgpjmB1d
NYuCCzTqpOM2VJH/NRpBPDHisKqjiwAgK0T2nQ9LJAFjSSlaEowQBD8ImNxtBAam4Enp9Mbg8eJK
+P/Heu+0ET5krawqrZVt6oY1YKlJiHMBP5PWd6xxZfAlt1KqQW5wJyemlHjasvrNiSkguZ0T4kvP
euoFBLgERK3s7eukWgdx4kcD3h1aWHURLmKdBMcIFpG8n7zEzod2kmB9HQKxPKuKJ5q4fr9WrnCw
IfHDk8TJdiKbAMOa2rTLyXaMNGmE41/bBoIS+7sF2WSBDSGsFgU7LIhZNixFw3N/oOLSGBkORh2H
L7XS/7hoivwXdQuhvyR/BucoJRZvMSi8Cml7Xw1JMo2e1AytXbxAKupOR+1YX2nuYScQDT/SF3Hw
6iofLnu6+ZB15WtNaUSzjkPmUt4zjKOsFfBhHCGkGx6BXGbc/G7kvxYTuaniwCNaDoKMlN4Ad87f
0fRAnwd+9uJbLVCZTORVujbfNEddQsYs4ZInHiWWBh52R6OXAT5UaMPRIBbtThfi9iuAn2upDH9k
nULcWHCce/Ke0rLiI/32ujB+gzSEXziDRVUhxJPhjBe7toAabDa+qHKI186vHBD25kt26y/TUiVW
YENVGBwee4lbCF8XuzmrFk87NnyZT8OrR1EAXHTQkKP75qqJ8IJrx6/T2Elh42nFa3XfY+tIqHIk
7frPQFQjuAk2Ej1gHcO6V3QHcuvbPC9WSck09OIxMqAZwSG6Ah1+P4ImZdQbsXaf3flDMV/Yvo/h
HGhXWCK189xoWpBuKyL4gMjtaXYE0zuDSbcO7dclLEVcKgYC0qc4Yje5Lrc4mAMhEpem0RY7tYi3
WMCAz9061Pb7Ew4kk+WMJqbkHPAeyODXX7g8B9TJV3ZMkcey9R7K9y0EzqOjchhFVzf0NIAxK9GQ
LJGqFqk8Ufo8EzPUJngFxhF5b53LvJqVYWdCKRDHLU13hf545e+Vb1MVGef+9WRI5E3+Q4B+I1kg
ACdGpcjwPGibj1h+KA7j26dOMLqq6ecYKRS7U9/vxBp9IXHcu/wvBZ4klPtiRdf/RikzrM3e4S0p
TL5IYbbqnZS2+IK6/2ThmdKzCqEnKYHn4gM2axn0L+3uhptXDRIIhpTP2otHyihAfL1URjeORh8C
B6XJpXsww/dgGlCtUIn9XvxoyGyUORLODIQ8ORSmHz8clrBlgMfOio5livDpZoTfMbHDlK6sw98Q
gGf4sZD9sNlN7A256LVfCi3mV/YjV90T0UTuBCgBolm2jOllb3oDaSUYkyIk9hPfqGhlFng73AdH
P8j2apGVnCSdh1c8Fl5ey7guR3synUbH4j1wE5CbV1YrZTAarBRDfgbvNSwPdUwDXEGlzKYIeqX4
DXnbI12S6fqWzWXH3S3508z0We9Q+E1L5s21PWgwQW1ntOeR0vCtU/AKvhv2Ao95qcwby7n1ZOAk
z7QAnWPljqd4H4PxprjhhUNaYnwHORJg598TBTI2yykjAQLFCUHgW5vgRYgVWsbJoG/zJJ5xbvTu
xDAVLfDXnp397UjU4fVElhjz9CjnidhWYqkKUHCxFjPUM3lRvGzeHf2pTRr4EASTVB6iGh0L9e92
daLGIsZa/eSroixP1d9k3nBsxYT2xli8VoknKNPhEVjhCtrEk+hs0gGeS9xlA6FN/o/vbp4XSGDJ
6IOumVzw8k0goR4f2wscOhc9sm2xl59D9TOLm+HsJfccHHSjYFxqNxzH3ZywqjLqTx3UK75ArnXz
yYwLLWyOtIws49LBq9qR7bNEp9ZX36b3Kow4NsjE7n3gOzVfRVwS08q+Vlttf53LRNkjep/D2IDj
U+JalwEGwWFfVU3dvms5jAWZxUDkAnx6Rz9jVk+LxGW3J6nrAVnqRE596vcZV+w7MxIyBJIHGsx3
AppX2yDP98P7F9XZX9FbVXQph3OlUK2O7iRa+Q+4NbMl0jQTRk7DOt658uOxx83tEK/SkTaEXYaO
QvRj+9Zpc8o4OqXD3CjMpYRcXmgRDCn6F0Mvaa9yVjmMKervoDB7ioDJWboX9O3pnmu78atzAxIC
7vMn6LtdFxXH6MSSNS/2WpB7O1FX7Yjd1AVtQ0BbNCx5gO0VQmWloH78+yWOAGjfpARBw+LsULfd
m1N+Ww9Ag9XAKkyfNecm2fyoEKkV1brXZaD9+fVAxysbrFg9MDSBfqSttdXlKsb7DrFwpDLxSOL6
/CPg+AwkOyKX1OmK4uR1+xqXdjgq5OIh4+Joh6VdWUo5+f4oHX3CNgH0mYN8FvglrpScgi9lVK9H
AibiixnNAHAqGX4IAAhimp42bJ7Q8AXp8INWghX8dhDKmgHUPK2c1TzZWYELikuc3uAVe/b3bf7q
3HZGckmDKffgBEuFbBYg3MWJzAMOJo4gsIyEc1BExZHJ0scS4rHShN4eXP/Xd18urosI7nH6fLXr
NR5N/Rax3Nhib8kNmLlbzh1poYQD7658N/PpYhPItmF7jtYVarTVPRjqdK+YYG1+ngs0txwmRax1
2mmcWVakq4L03qFtxoPXvyHcnoPy1eSycgahkKAt+fds21AF3aKnLzJ/i6Vt8hfZcuOPUd28Ex3K
Ak3iO5tyoBKC4SKykqC7n4QXsRiBO99GCYvLmkCGf7BSt43Zc/onsbQdbJjI/73zJVRz8ElAZMEE
qmS2c9gz2M2fyoI1e8tY6KZcMyYhMe6hI8QcH6rBim8ryAuo/45wLkkCrhVQGrx5ARAvDv2qbYXN
1iefxiy5Ge70cBbL5bLIpfoGYBoHx4Bbgvn32hO71FTTMWcFiZe1vhrQZyDbKKKYxi/ksWGJ7YCB
h/4uIgheAk95E49AVKAIz1YCzcryPzt6en/ygHjYaD5Ouh5l/5KJYso5+rd86Jcw6KlA51SlwhiZ
X81Cw4tFeHkplcbN15E1yHgOdQOB4sGySf9YxbO+g/bVcXZFSiqUH5fnTYHzbuiwjhQKaseU/pC2
XpAs8mSq7ENVoKKv5K1DHw3bGojO+qKrTuXOZqD6S1U/RuTWhZZPM2qFZVn79wDbWnCVNVcQC4me
AabOjaN5yl6dxeQa8PRaCP9vNhYXI9EyUnkH/yerjrs5BQ5tcm+JB9I2nW5yLbO9/d/l2Hx3t+ei
ROkShJr7jJQog2mOZCJrNCWnSrFsdtqvFVvYLrcz8e1o4daGsTQw+dUHyA5RQD3f4aZZIYU6blIT
rxRkD++K5WNuN4gocAgLmmrrYPpcC8xKvO+fg5+1SW2NQsTwMSE2v7BQeUntyQYsfTJIQ8qDz1nF
YNRbYaG75JhCQj266M4Ail8vOF8+WYNZuOew06vvExyV9PI1DefV8CQ4R3rI75ahzXEW+gsXzue3
Sp3wmWA+KtLSg4qZyyjaGIITV5miiw2GOnXcO2f6IyeXZdPG+CqRvShLW6ejMrRzYtqyflsQVgnw
P8El01zD0j/jUja7Di1AZJIBDtpdSU5dozOnPUXmTirSST23m6gNhuIAHtB9L3R4aKyeSy2KIYvz
1XhEt2XzcpvGD6fZVnoNd7JC67by+GSqx1N49aJpE0BNerU4ZEVqM0Zt7SWX0Z9gTY2kTAM3eA9t
lwT+Nm2SH7nR9pZRJXS3AuvCcQaDWEsd1GqkEK88dU6PTK4GTvjk8q+DMAcJYBuP4nilWnkktzdS
pEqOOkUKUueJDMFyFIArBrnL1JahXMbfmpSDJZR2BkW+GvtzWP+lAENuacxQJn+IwQK5TmKKVNd6
9FJpKoGxwnJ/KdDZWL3JzSlKUHyf30TXdNPl5cmGynZG56QdgnKQZHFZ0N4+l4T9sWMxNFKPOlAv
knlWsNNLlwvlSTMiRc/5KM21QtWr9Q3g5Hbrd65jGtDXQ9gud3r6eg1Yxnm2A65RSnYE6m9DJ92n
T21QYTt+ijpTqyk3X8CGryiZinKzmCVXtcYr43lmKhNHBzzi8iDzNHwktVYjLM18oRyMNp9uVIM8
akH8tgGTUF8mS8Yrlr02Q+mAGBUPam3R3Gi925PW4mYYsLvmz/B+XHID2ybrGlbop1oXDfmNz08d
kCyLOyRwUxo17Ve4HzAGz0S2pFhIuYov47Gxu0mDjEYrlCPRlaQ/qqXI1DNXpyqZy05SwAD+2smv
43nsCUrrTb5ijd34hsg76OWbEDk+VTapjIzeM1bJdHXzCszEnLT2FfqYeHStlv9p6KpZWthd9WmR
xtvjtXcxZEdQxyfRV8eriYRIaINCEthzsN871ZCbyDV/Ps0TA/eK+7AiFtSVuGzY77UAbl6vwNlM
TCGdy1LlVv6tSMOBYjmpk8S6ehx0i2khXHYVlI3HhgRUv5VLqOEEg4AftkWBfTeOR2I1ZdJEbwoN
nQf2NzS7S+H0nNdHDUeKEiZuUR3vX34hW7FaPIYq25yejBoXBV7sPrqcTKR4aL/Pp5Y1p7M7jqoL
2bSCvX9G7GBBkwdyNzjafWN7QEh/m0xKoWJ0CQQGNFOCQLjeCDaJtomOTFb+K1vgSZFsWytkWH5K
qo9X8GD1mUKIoS9UoukpRHNe7n+bd9e9hmZJCMXNgBKFhO/9nwIH+LUzGNaFNV+kGxs1m6AxKzVy
UVr2LK2lUEH6OfKO+97N2FjjKwgK5e78WwozxjtHRuuktgrrcQaGpy94qjDf5mlEoFEZbSdT3ISf
k9UG03O8Dy4X5jeQX9EGId7trx1AOyDoiOBqln7HsXPt3e8AXSX51A9OX6KYrNSX7EomsO9aobaK
xia5Rk17FRDIkcRxFvHgQ65ewa7YdNvaro0D7bTWlLar9ZjOD0HWUKcHDx4MAecUBQhHTtAjUvlU
b0kt5zuCnxbHY76A2kxAEyuWclIZmT0W3eGNfvdpy57iDFZ2g/XZhgADCnH9NDuJGTpJ1i1ZpF1N
oFZHm4N1RqFOnzU+dehRInNDXoH1ns5De8rlr4YWfx/jaxpW7qsbdpsdbnHSg7qTAQtkl013bdZc
ls3lzwCp0GFp/4pHkZaJ20WW2a/jTOYeTOXOWGZ+yCHd9TvOIse6xUcCpbGmoh3nkhPOZAEDhFa7
pGt3VtiebOpmYXD+fJmYcYsMFwMOT5pbrFJKyU7PAfI+bR7rtTp73bgkRsPniG1nx14tZPk3BoQB
lKm1xLW+7MAi0jx3swzcRWNWhgcSdC0guo1BR3Eoz7Y+ud/K9tdaOEhG5W3ac/q857VpAjEheOB5
Pi5mo5ml2pQNu1KgvfXcDBdseoTpQmm86wFF3ILr0CXMADWnzEu59xi/LdwFs23cWXOmdIqZZtbi
JMV0pdVmp3C66VZFgBzSUcfzOxSUdk+EigsMB+Bcs3aeyMluMqu4tay+HMY8lpTqQM1oYn6uxZIy
/5jFZ36rihxPPWWEseyI7rtJFr3wIErT89M9HywNdhDXDJvPWcmIFdeq5QiJg+WH2+/taw4yNoTD
UpkZWjtdjXGmEnmphvHfDtZaTONowsSWnyfAMHR/vFILt0GGb3FBlwYlAQ1r7ea55/MPpiMWMg1G
n06WYdHFRQQoMHaYOfAkd5uSFk43o9b+w3Bheh0PeLWy5BTKVoO7VaJukptA1gQgUnNMadxxe1No
rwQvzg4gcc+QYQCaFL9xNBgyMvsiaYIDc0Ido0Lw3+ZyGXYNGldGndqluaKyhVj1aPsYO5kT/qj8
aWy1iw35CKWWq/K1TbhQYvWCyT33DVElLcvmhFLVZBuZAteCqeo5PoNWImZLY/d2noxhd0FBKZwh
6Mu8p10H/pIIIcb6Rd4aJutjyPfr604nbpJD31lIJ/KS0zVwUlJ6AbDSdou0uTYyCFJdaSDYGK1J
vljllMK8qWRccXib9SPCng8QeBddRHOTo6euXOEkvvMYSjjMqQ/9zbcPBPESqLVzbxBbHW/N11YH
S8PZXV+1p0BM2R9jghQWPT2SgKbFHrP+9uK0r/e1b639zDKKp2GRmQhjGhScGvjq4BRNhtt2IgQA
cmQfIJnwfm1giZSGaZznzr//oVYFyq1IaBvb2Lbs117z0i0BPcPiug+Evo+SQKbV2Zo9hWC8JjsP
XSMKoVcwr2j/nSJvhGuHO+WnqJZ04zRx8Qe35fIjcFO2mGITp4tHB/Teb42In7/8SXKjvtB76HWA
CS8bOMCjQbcyD2hNUK70Lw/TvqhFPKYZ7c9H/b3EXs9EAot67BQ0aoRF9BgtHymmhAoy1KAalRMH
PC5S7Xpnwbx7E9z5DWF/xCJgoIUgWpb47s4zD9ahZorAHU27mb6C4erq7HXamfwZCkGQxZ3zgFcM
fmI5gz4krXBjntyefJQ8/gsfujwnnGUzLR4r/Kp36yZ1XgO84RpCZBMwJqrek9sVYjEjgqt3lNfN
X81V5uv98b65bZOGb621fqLxlpv8CqgR4d2KFdlvgosw1jrceCYDrW/bD6ROChYdY7Yzmu6zoon+
yNAdqLd/aM08+G+lQTnEeRPsGMjIj1Zx2Nhj3wqMMfjFQXPWztNsCL3BSqxgBzeXKPpcIUjEA/cI
6CL0Z9g8V39s0NOAcmmdlq7pKNUMFO18nCEi5Z6/5BZQUgezwAu+gAcEiPVfb+oTC3lxW2XY7jF7
Ksfxdhlv6iTbd5LGtxZWkeIBcHxTi6IA6uwmmRoAnh1VWA5jd2FX/t6WEA9bm9iqOL7fpk4PpIWv
TUA4E/GhYFFIe+0ND32Nh/1XWju7as/tNf7xhqFT+6HiJ+zpkOnCOazICtX/Vy6lKrTEx68Smg5T
dP1mCxKz0ZQzwsXyeM3r6QOYx0hI1fqyaEcsKAey9xuIgEnJg7wtMsksNzMoWiunIIfCp5fQjhLM
2xhvelchow1o4jQSyUzJwPsDjzm+u1b/Mkpbfgz0SgcOoFYWS0Btgn4B9sOI4VNb3taGvRZfWNvb
CQvqbhxxspBrzGb9cYd5etM0wY+enBF9XGsH2FRQkIOZ5LhRT78+UD/ozP1Fi9TE+memaBAktp5g
JnuOtVRfBnxkicst4mVzTPVKMc0Y6tPV5G+foPSelRm+/FUMHdncIU6iQPk9hvFDMonlc7quuqsL
/PW5g5aMlqUH8gm69fXnEswlHm0mALjnz7q8LJDZYjbDaPzDbVnTGEqHSePrk1sB43shvO6PVFN7
whmY66o6dc3bgNEs+rMUkseD1IHneUWf3IIowTc29Xv0zW1RGIWXH+nHsn/i9fvCNjFWAeLdfmdW
kE524lKyygI8/FS9+HauWSt5et0F25I7zi+Rmdv5jEFul1/8R8TKYKoM+Pjh0mtGLYxw7sf1HD9L
oedYaM2v2FVBZ46CTR1L1u8Vd7uVBsMTsTKlHHsNtvpCXMn2c+osK7xKVGrsL2uCF7lRuYguz5h8
GFY4pN5GYfzPoy9qTfEqx8/fXz33tGfLa878R207M0k0s1nUvxxdzdDewx4QqwnJjEqexu3rBVrd
QEEDsy8dota6TYhf0Ef4MhBH+pI7CygIQ0RHefhfimZXr5aXyKODtA79YDJRnfEXZuGZgjK+HjWm
QZu14qYOwlsEy/xlKTqRmlMWcOGmva+mKlGRZDce4UFYROdofeNXtXL3ycxNz7lYNSLr4gBo8YjZ
hABhi7qJwJVMrS3NtRLlLl408XEVCgW7NbC/dAgvrLrOgwz1WKXV/KO9QfdHGp8j9Hc+ZSr50Ljr
FgoHmM+ZPX35XRabzt/sg00APSVeJpx3IHS+2KGrl5c/V6FZpfCx+mDpJmGtsATPbAmKXAUavJzM
3IMTmpiWPXK9OAXJ57YpIQd37fGu/UNZ2l6D7o76T7s2GKvC9hO3AQYlCiO4ZtrxJ3iSXF+U38rV
8ZabFNkXpPnfhR5A0ms5UM/+hGt2WGXowJ4XZ4vVTkP5TmfsvtKxANot29434RgsT+8COR8VewUZ
jq9JLQqBrpkuVWkkIwmnFyrxPzuY0lebltPMxUDxrI+iWI7IH+fBnLKx3ga6JEOZpW2Au52EdzLb
GB24MFmQ/BDxd1BwN8IL3iUUkT1GPY0m1efrPfO4J1PbV68f6SY4FfIdrJb2OQm/LYRWFSquLKgG
R7vSMA8CpFkpw1hBN97Hv7MoS2d0126s83f0IDjaVRL7lNYf+LukFtGDOKpYIHU+PvyeZPZDknm4
o55M7qMXckig3j3re0uMKrUQlteH0QCoXiwDWbSIvAbyTVj97kdEgYt8U/3jA6SqSyyU1qzQz6/K
W9jvfyX5xm+YU5kydxseAF9ZnKupLo7F8umVz5l4jzkrQhLi92uXNqMWR83n31C/5MxUaKSnmkDB
IfRFMY061UtzjxIiNfnBq7h72hohnSqz/V+AfAROcrFIzHqdBRMZW2D7glhAvdSVSBfFTn1bLX9p
rw0gCyoJjimkVtPLQg/N85c7O2mhnSAABD1FT3qnh6dbEEwZG4AijK8QifITX0osaDZSGTOpkKBB
iOZUQh1cxqH0DgTNdJIT5Wjm47a7XTdgV7Ot65XyEKAi0XIPXMFvPWRCO411ppO2NoglR2p+LIVC
rrVXH6X7fSbXzvw3+arxVW5q5GwHqARXtE+vcag3EIPp6MB5tPScK1tRNj9SiPfE+Li2xUcF/gY2
K2BVOkSVLyhWYLmx1bbs5E6mne9doQ246nsR1IXbJinPojiD03v4wQriFMY2Gz333nE9hgs4b1ex
kOd6LVJJSnYC7ggMHL2SSfn6ni4qJ1uXcFQiTUlbkcCZKh/zxaNwcGdkc6YrlFvnQRxbciadoGpJ
UBsFITr2tPH5xTTY+D6XUY3mqmR+5zTWhUEP7Uao0/57MwgCClXx4vKh3necErU455MOK3PDYsUo
KvTfFQ0p5Y6HzKMoMWPl84fQW9x/PfMEcZ3L5sPE8bUvmNko8ketQAXWGKdkEdhCychMhvc4YHUt
uhLjrAY2Lt82sWJGc/NUlyoL3El4rb98ilunOQoOAiXlFMS36jpRATAz/tbTDBNRpBQFf96uWV1a
JnFVycUct0QogZmVzmeaVoNyOy22UulSSGalCWc2VIsedEM7Gs7/z8uthVNGBbBX/KjafaIHgVkb
+0dnaXC1ef9DxAtHeOjwrN+tFgWNoSVY4V7EuWI7gr7I04tAbQ64iov3dDqEz5VZM8ka4mJdiyaD
q4qkzjVxNq+wh2Y613E9sxpqj3xzlvb9OXONJWm70m4uzvYQg0g4LHyFyOOCbOalLBpxSAkJpqiQ
XZYSybBuPcTp/a1MFiJgT+BpQ5InelR4K1TWO9e7KpN6L2Xf1xYeKbGvHy9NfXlsEpneLRhkey8j
XrYj97TMqa2Gijj+is7wizrNgx4LDiXppZ+eYRkdL80mqMdD7Ati4bf8GF3y2zXYXtuAheAChVGK
8driQYUIr43Wnme0SH4coH6udjGZuof61vSvHNvORK/Q7WcUPnCqqfCyc8Qq5OLLcomQfFpKKM3H
34YB3l18+9QBh5i5X3C+TSVpT0/jzqUklAyvKvLJoZ6x9h9hrsHNP71jZ6z3bSCnuggAuPGogofp
TY5kDYTemJdue66duv+lphE9xK1pXAEuyaHDv9ScUVXesYXH+D1Izy+hUO6P3S/FTY44LnNa81iu
auDdV+Np8hdjAYLiggfJBlD4ngP8JD6ZmZ3249bzR5Y9dvfd9tJpb5b8UoP+GFN3hNsTqyOIrpOo
LdLBjRyhvLa0zA75h662qpZhfNn2Q5qdqWrLkRammsSrrH7/0sqhr9fn3qMxIXP9GwKCsNn3q/uo
2zAywc6w1g6sMRO3Er7yH/36YDoRpbRfrarN3C/0FiDFKtmi4ijgMObqTHCl2eYItZ2JvC8+MSAH
+2TPAsLS4+NOFudx2ltQxtJGD8w49T+lTM2t8JRRzarDhjqAcxFrgGIN2rig86ERki43VrczTClM
iTqteaTDwQAVGycqWt8imSSxELtsLCyEYrX21cbmP3OIL+u76DUl8lX47VHlvAJoY2kAPOayaBRe
ylFGVa5rrdRTAiej1J3VfH0/56QAsCZEI+Kc3sPHCvAdGEdcnxpQIHpSkULqc3HxJooI4y2C7u9c
pDHoTB59IvTgyWXsFrUsfsOjTmPy7YG6szgMcoCrHEpZE2DecQv1jiXiMT0bEa8wDE+q+fluskd7
XN5AiIn0/5DLKyEvfI3e3jxJVZbLfWig4qBdTgYX3CG7RYzfYh4fJwmoH+sTkDtZUJfKv45WWDvu
lyvZ9217p1Up6Pnp1aCFV1LzRdaPAuCRLwGFaXhX/YHpiXZO5UnQsrpyKpOacGWDKx7iZo2qyGBg
s2v7vIGR+W5ln7EnKwLC7r3vCzRX9AWg1jt9NXQtrNbUhWv99cTV5qdPXSrJxsqxlbcV1a1AWDUA
yhe9Uzd97bMVHtdnSu6mMaaxYUOVYRBdCgoo531uC7hJchS6BMYAcp+iH8cnF+rqTHk+SZOWHPzY
UMBLs76TvPIztVD/frvMH/iN79Crv/IKD6qnATaTEpZTeqcY9YlbYvPNc9OC0NTsqFJFKHE6E4Fk
pCs+x3eyJTYxcr/+pIPhX6+chwD0nPH8A066kfzUoeDrrzfjkEDDQzhRgVbLLjdKOSFkDAm910FP
2HCL/Dt3Y5G9oIKk63t/Kp1fLAAfCMN41WDzuWZiAwrXglEDtt1GykIRvolLNq7xYLT6lYcSB+/F
2cHiJVL85TsacZsKtKT7yRMSSPjEh6+lmONROTHif160o9N5SySUzHfqVpkZrVg0DruWx8XCgCkQ
1FMgzLAYhgpklquL7ZbnEhXz6QNAiogDIAw7lmdAPyNfuIu6m3FEs/oraYpmVCYPMusRdKSieeHL
NYEwnAbtwBDvn9j/eWjHZYz6W8CkzfIHxkZfYunUnUI7Skl0OsEo9KJjmslFVhNh9Gy7e2xqfNCI
ckXJCet3b8yr/IILGHZG97Q/3QDBC6ICH86Fo6aTSOmApoYoWlvGjR8VRHzC5GqFWVfvpFnvY7Di
d3IUArGEs6EnqkYlDzMQLhfBmjvVh2CG2F2CNjIvm+4u2DikXk+fV58ePrZ0zkOCwonQWLj06XCi
xsTE0XXvdRFpQ/4c7+vMM1mJcxooHfrgRT/CTDbQOaM+b7mfnTz/Z0iVR3cXsal/XcUXDGu/8o4E
u2w+5prFqbjF9bXxI5cLudbUGVJlDXGTW1QWiDIj11hY5P4N/VYKZrz0yBopQ5vQy3CsEP7Do7hD
g8TfIaHD8rLdRID7oMi0C8LA6d9Pnc1bksSO4WckfubDMoFEI62hBRyzIlV2wRPN+QPPi81OPBq6
583ZVWRqYNDhzrAoDddfw2I9oOrJfsaGXzc+LmhDQGQT9js2mzkUOyYwneoBTwItXYE9CR2MsalH
QEz7uV/i+s8ZLBQOrg6qtXXruSc1DuHsFBtGSO3UvBZHFJjHowdyHRhYlLgHKU1BD1eA+hjERRPZ
DwqeQxgwlhs/At9ID5Alo2ZqY3YluoMcPv57wKkG4uVGekXIgnbhJBSu9uswDvNS8NtEGxXPNEhF
YVrsTv2SPV/lTyvdLgTF469G/vLEGPh0mPZ2F9u3a36jSBRQgsu5I+i5gYN7lU70gd4YgE6v8DtV
C5xqksoEwK73sJLh9DArG9geftEcDd8ojB+ctfE48Og0ZTRI/U5VtibuGHl+G5NKwuT3AGAFrBpJ
BK7i9q5TWE0SzsA++PhjDVc09IAeJYho3qM2JwifU7p0WhR46mNLsLribCfvj8n1W/RAJ9meuTHD
FM3PHuw129lUWjhCPjV2mgVnixR6QWWAhIaSkQuRgCjCQJbVEhqiXDe/0SgYdV3i4397nTaWMiVw
m20qqhbsSHVnO+SnnqL0Pfmi/cE04OzVZZmmMcXmuAyeI8gDN0IxfePVNpqj2AbxQuUoR1Zj6uar
Wpfgo1XMZJE0byv5SiWK8Vec4MQLBrKC5iJsVhwLB6Lx7ggoxMGQZxt2NffZHaIT6m9lL2WALJgT
cluKSYjt8zQdMDCFkIzlrDFkwcQ1oP8To7/fNDk9uAJarQ7h/FgBbZF+exVrGSM2pRJOoSDBq5Va
xSKozjVdvSusRUhuAqmmGqF44Uq1UlWC7mmz0IJGkwLYSoH7SF+0cieyh1EIZBCgv93PZPsVQbBU
rcgpeoglUfKUUSCfj/KUOxyfKzBs1F0p0j0HABjWOnMd+i+JZ6upYTStTgy5l1cymCKvdX1HYwtJ
gwsfsgS5TNB2jdbumYiUSvtWDpReuutztTk4PO+CaykH5bUmZc13w/iIt1AlAASUKkgzGd1vun2t
sWWjRtGcpYIrXai/4RAUUCHH/wa0/377VoEJ1Di+/KBKcYUfc0RIjXc/wOW4gQY/0cvRQnvc4/Wb
FrAKehT0mZOUAGfhUtRVkkxVnOUPHEPSsXkAn6xw8dlzr6/rHUCZ47cPgSPzx+QFT258uz1bq51g
7B0TmdhX8BmIvNoF0POr93EV0ppOC6IgmnRoG56mHCVOsIHU9IIvb77tIxykmqJzjvLECAiNwrnQ
xo4RW3WpRLXogRa7MdN2W02UndfbPYJaX/GderftwRhDjHNPphvGSmZp+PA78g+ClvzUsWcvrxE1
TINJitP2kioMBte4hqj6qBBtNurJl9Pek1vN8LVUCoVja4FeOxQ8CM5AyZ0Hk7tOC/HMA4qlTOua
kqlBQg4lxpqaEWvQ+HUefuivf8C89K48lnw4nO8bq0uLSjMs/6c6hGpcLFGGCU2GZQTc14X3RXbW
988mpzPI5hckWtiLEzBGYzYhBSSo5HYOuoxx4AaVmQLml50pdY8GDtJk9+nGfKe/E/ug2fGaJOpR
6YHbBATftkoycMB3LT+JjNZrR3dgiv2yHU+zELAPz8GKMFNRuhk1KE8ay5jFRiCz7li3pONfj/WT
Hb5ySddVpQ/HOS/RYCq1DIs/9KPsc3BvF5pp6HyLmK77TC4ZJ/m384+UJLWgoQ7TMAjyEvkAarss
diJjIqn5tAF/ELAbcbVHuSgTD3fyNZfq7T9PGSjq7vLkSNBUGpQDfz4aW87JwFLv854BTkT1Pil+
gwzppTPav1D+xCT4LpfGhrzXlw33ODqin1Zy9VeOcGhc1qY/hVD0wPYVFR1AtUOI+VIrFzByML2O
DI6icRqCf6dA1yUd8leqJ2bvwiTPVhad5a8G0lDxZ8cMwA5AbVC7FHV1glVDwSy+SDaWRs+eVl5m
66lFlf9jAMjGKgNgN4d04x7YC9ha6UIQfrHP6l2F7IlnaYiDWcFlaVYbOaZyQwY7F5M4ngoRt65J
WpFJZVKP3/BooUtc37biCi+qOyD3kCwN4KW2hBopgdwR4P5H7/tWYDjgMmd+tKG1A4vVv4bUPJnx
jBsdkI8bjzJhTKtxSBEtmx92iMjhUKpg/LlWoNNFpwBkWUrMc30iS4YTBuUOIkgAkx5q4QdK+m52
NHtywkPW76jv5VERdDvFnN6JZE08l+//McvhRVjPyww0yAMLbRuHaqQsUWnzBW/3FavYQrNL+rPi
cSViJpKobpy77Fi3MKsDkQ8543tD01rf5a/DU/XLOTpSN5Ndg5aysnY6hQw+l4XygUei0ieANEEQ
xaerxKkRw2YTnwzdvVWMLhDmdWcwCz5LOO2nEQ9QMPfu+GsGse3b970GlKB7mt/9jQRkNn2VHU02
b7Mfu3uPnwWvdl5fyCzbQ6hMiKJGC+fTloIu6037fdHHtQeaOIgWcHkCQIj1pmFFa+mPzIukFuNS
F88iHGuoxa8WYu01OOFJ4c/K6mcIPM0ASbYmMjvjaGg7L5/EWYbtr0skH8XH30DSzxFCU8wQpfv1
FbfLmaOQIOiY6p01eWkeQYoG/PJRUIxqM7ustw5npPwfZJEXnqQPziSxFhT6zgkh9r+FesFAuivX
mZFHBi6nU+JJVXnM8ossVXX2Oi48Z2Xab3PeM9Yo1WyyaFb7674FlFx+Xla4EMRVSm6LacE+ZqFj
obY4a6tnrQkAQn4eZIT9k9dg+6OdNydGarST1LByJURHuQbfQmXPpiMQt80TAQkDm0YkNx7mxlbV
O1cxQiMOVjcQ9KIFll8dtd8dMZHyG8CGLOQH/ydy1rWZc5kVT/ReuEq0V6WGZg5zi5DzzBRLf1Kl
fchzkHGXSPyzWhV96x6Q968YLZsNstJ0VGzul42hNVRj097DVjHgJ8JBlXlNIFnUrvq/TFRoPsuv
htEoBX9pgvJzviYS/K7SMZCalO1okOfmD/xwV7zgPNtJqQIznxQqJpoy5o6YKMDsK6mMC8Ad1tFL
G3n5GcwHwbgUoo8S+w8W7vuJ9c8MCC29l0e+UGNW8CjC1wTukAduYn8Gv88JQCwuz42BdTDEmyiY
AdYZWStV25s/OHuMJxTZ3Etakyt4WlN4MtLWewrvovHTHWs2ufvSVhAie+hjTf4Sq77a3ZWpA/8C
f4R9oPtE4ygWmFJ7jGLDUz8FK6XSrR5LMo4P25cs3vURfITc2o2xQbJrH1X1q6W2sK4mTNd+26wl
671Hc4HmxywqeD3BQsrNYXKcBQvjgaEgxn3Krb37OvQTg7liPvJoa/9zDur36kK8IgGLLCbG56nJ
U62BFS1LFQGRxWXaMTEXSz3fm94BnSMNLL7lQfn/LpVAl0ajF2qRqbdwqaOP/x72lG0mpG96EcDB
lP7mbzWtCVbO350vdEmfdUHe7CFBzRs6BIqzDLIGSxVurX5iG1ebPvCReXgU7D9CtXQPuNShE6Od
wi0gqCf6DkvUm1CrAPz57jUtM+pzoUrljyjjkAsJDKhFTcM/Y77jNuymI5wflL53geDdJJHiOE94
AN0GgMe+gG7j2euoViiJBryIw4LhAemTP6ZKNFP6xPAz+7JCFDCIR9H8OPQ7S8JbxI8q+DruWHr2
ufqIfhWfrkjRgGdc4EG6rlT5QBdo0kRJkVtd4KChgtfCpHXvEk1aE9o+SssDxWds7kee/TyG++9q
AKjd9BIcDk6f6uajAMSt35Yg2js9WVjOlqEA910yVyowAzCFADHvxhyZ8wPDN8AWQe/fkRQHE9xt
uuiuWOlS1Mei5jRwrUIMZ+ZnN1YhKd1qGeq7rH0p7UHty2TiPY15qZoExUkswpPzvJGjowIrcoZq
WkprED2SGYxtlgRjSm9bwd9zwPZIWWRH0im+5Oa69pWKA+5ipW3M0RCl84AMSorszayz68y6GM3D
tsfnSayqPKUHj7QzsL5/kSn+1z7UivPzqncE+tVzejO3Vjf8M8RUq8I1EKjVMK+5REBq179N4fEq
zgRz5svh1kY6tO/7t/91tDg3KLKEw8Hv0S8QOYiaJv/aKH+/P2nJsdqbE/M/N3VfbdmFyE4uGKAW
hu5Za3PqvQd7OMlx7e4TLWpSg+OgTKHnszxRcNSI/g9gcOLykccIz29jW1U62Q5TPLmmRgxXTFY/
HVspJvRPIk5iRFU4YT89xz/Iw494CUye6N6UttucC9EBNSt6bsA9mL4xbsk7X3IntwwY7U8+CpDX
jkBBtAtEg0e5/uW74Uio6wxU3G4Tueg7GxQT8WDAiikxEk85n+DkPawAAr/fBLXbbJJDUCk8GjGI
GZXP9PPvwXwgX3R/I3siIfnkQS3QTtRY86OenoUOtv39DA0KoO6JU4efEqYkgsKPSvaGqQdg+bGr
ylf5JS8wjLtMKM/f+oIa9tfiG3BBbnT9mm0Ef7VNuvX2y2ItNR+4qxmeJU2JhqGo7Gg1mlexM/3F
kEOIt3qztyrCYLrENb4riH6iBM6AUqqAhkjHrvrC35Xr39gIMn+FoNW669VQAm6BdRrHTJVwivQl
ZpB9bARLVgWQo7lRAHpgu4VL70iKa/Ljv+KNyLfmXzWGMGJAbj5NsQVdNbr0KoCbZe/oYyHd7wdO
CVwYhGiwLSfWvRV3RxS0NMvVkG26SsBMh81jnelsHH7uNlRh+Ns4/2oyzzazYywfL15mXEcUZyH+
QYaI+qbJAAO0VoKWWBva4pIrp2OgSw8+s373JSECF9Bp79mco+AjiiSSjdTycB7VBAFW12pAGdcm
uUEJhslyq2IzbHkmNDnqv2tlqBFIFoZjCBkjtIrzTupeqqccv+DGwnfCTljv1OSc3/J6WmMTAjdb
a4/NDOoNZX9V7pqF/dl9zV/tHj2utg7ggIDUKmnqTHHb/27xICYLMiM5/XAfwHH0BD2vnmmyYlD+
dLqJMFnr3PqJCywNl7kr7lT0ruBjYZgzXs6ZvMlQgCwxivOJTKS8d0FSMnkx7QchMeXQ9IwWBfZQ
+jBXlSI1Sc0XMENycWj0hmstSy2+NM96PGL/NTew159y5dYGOL7Bp/OtFezjV1tSxYOYbHUlJIAl
A1AIQvZNy8uZkap1m3SH3ZRr87EC4CGxYZOZ8CgPmumT3NIdLcTlGJbDAYh4ooQmX7xiLnjRIDnP
tuVFRljB0OyP4d77RAXJzUgUbnuDHnr9nQEGNgUhtQlZfXE/KvoJEqyRkG1uQP5DbfXLG5SUAfRd
RZMEebkd/X0heFahFdb3ZUa32ItDn1d1/pbKbZWm2ErXquhYQhdhfXf8VzwF1ndR4uGIeN4AqPBh
7Oz0WVyQoQ/UGlwSadX2h96N/hRBsaV7O2WcIrTGay49zcNy3zM7V4j8vXZGD6Ga8cQbd0nckfWW
9jebE1+U5ygpMqzszaL4Ahq/ES8MNbGGy0PoPb4CEcRGFZaOnTO4jHL579lSeJBtY3HIamAg8gUH
FHbCkga+MacMQPI+d7OdDTf2LgvMDia9v9vrVyPFzgphvW38Qq2evWiXHGHdnnxNbyQ23Dy/kYdy
tZvOCImkL3IwFuDsscVNjgXOdPLFPxxKGlVqKfHxWSUt+fJZAPWEDu+38ZgRVdVqi2rlOUtWJ90c
U+2g8xJeJgS9nKIAUPH873t/LPK36gRdG31EpOFW1eT7FZLpPsEL3uGdL2eHhBqHxKIv16s4JLV1
GCUZ7S7FHmbKwULHZqy/DeI9jxVr3Y2a2cWjUiYXKdbExHifWGb/A3le0aW1TskhV+p8erUFfAt2
JCJ9J+GFQdJS9T7CQnOULcJiM8fslG3Ew7UF22PqVyEAwQoXQqCc8IxfwmTwrYgeVrexv/oYxLxS
8hW6oxbd3FZ+iNX0DqBW4ABQNcMt981EBteluzP9lpfygTXN8D14MBpAp1211H2dpqdW551nDL0y
1WMqL4+3psZwTPtyQzTuZNbPCaqYDtXHQxKoMtxos29yWe0rZNkj5vf+Vij90QZS+sXMB4xLhq8A
HHV/IRpSALRz/0M4Up6T1jtENBM5s1uSI3lbM6qEf50nBUiveEFykRQLLrq/AqHEvqty1MnG0m99
e/qsozbI7XScy2vhg/6dMb7NVAUb044mG0Dnwz6pAnmdwgTlW0BPXJ79mULqHmEkVw9cAviHku7q
sAZ5SrAg21GnqC3QdI+HaOyPYY5xE6zDa2TDzto2rg6fL2A8chrWBt6XWRoXmyr6LkDxwKgndIsy
IOG4PvRRGhqru5WwpBXAsEI007o/2zIzfYr/biIJa1+sej5SEPj+81NDDilpqLc3LEqWByWyGTC4
ufQhXiG/jFRRoG97ipNDMglEU7v2CeGGrPYVW7U3HA+s/ErucHjEmo++WjcYYYG7h3qKJ+G6d3So
8RFXPx3drbAlzC/hJJ6jrXWnPWWUNN6azO9fdAoHsJT1d3A+SClTqEj5U5AkGy0TmHH3HZcwO/JR
2jYUnGYxy66abjPZGFTOxgAZBNahJMAcZhSuZsGj5VghHYxlPu38s+I+50Iw0iGx51hNmJpjzekw
mDltPzOKBHJ70xCfaWjVnc63BeMJaCVPLkdqwhmVyARTSCAyPpWfz0N8T++0zmDYFqn+vs4CaKfQ
c7NgqbyVffy4P4JFbB4VXGMbfdTq0C6qd2GkRPn+96Zdmpj9kTaDET938B2FB34596iylRJVo6bu
gMy5PMJQS3e9bEBGElevWu3A7Msn8jy2ZfIYr3kx6Vt/b07wgHbEor4dnEBod2C7rTpbR1cI1Cot
MchRqLSab7I45HXwq1d6H64X7wHWvLtfgMAPGI5SXHHHPK0puTtx6ROs0kRlA0UFELWEZyPm57fQ
sQQi4lhemi5OEpYNE3TwPhql0mIMwMZAGd36B7z5/eILekaw9KSnP0Q9YQ5zw1oxj4n0PXgGg/Z0
dHKUQb25h4uDzdQoaIvapN0DghMZGqNe1OAAHlZH9RsBmsc44xpPQFxaGNmHx6r4L7WDzxSb0V8q
NafR5KjPXhU0lkigp9GuvVgKbuCNTKfi+u40Bms1iUdoVJPzusZrsmMjciQkAsgaj9Eco6O+Vq0v
jJ7ditNH4RZmc9ZiLVL8GJS3HQNk8ov25Otf+ZdoqMlrCAuo/Yl4xJU+pYiiSpz6DHKO/DC0EN+5
etvCsfw/kQxf2v6mX2ug2lTYAR5JAAaQjZ1Dwuq14XRlCPxqbAuRoBz4PhixFUv7Ejo6Mcd8QdQC
3DIKjtWpRMy2sx+j1tzySF/UnsdWRDRsA91Q39y6E7gPj2bNwi5w4vb8DG7FiUDD+31N2KOF0djL
FWbLlbfJdL8aru/jGbC/NfUhv4IQhTB0FffRvhWZdOgW95EngEPyflEFrEXLICnmw/LC8Y+KriLX
6Dfg35ymbncgS1pD/TggCtYzrrdw1JqtaGideGSCofQsRzBkHSqXE2UIaptNMphtzruXyaWbUlmz
wMllD2PP2bDY7sNgBifZbcrpIsKNS/E13VAW8AE4wYb7cxyPdAoNl9jL36I2RONR1X+v8c4rQvk4
8GyiLQJD28UfeiaNxyg6zcD2cv1RjDO/IA3X5JH9PX5XrUw+0JpekJZ2OSkX6N9xBl7U/sNHQQy/
BaDzXCHOf9pwZuHY8l+b4d63INsZEziPgHnTu3LgTxuyFLny9kca1Kz2/yy8yGUTED1a/i9MwQtL
r7lSqTxYxygqhXVhBXu3I8533KxYM+m9z0Y2igst8Ack1apEleBfZ4otJTCHDrSjj/nyYrtiAgnG
vHpF6R6I9iTstMn6j9f7YFrsZ8m0A+bRSEwSb1YlFCqsBTZ8gH0cyNxvbrGpw6Vc9AruujY+OPbq
Wf3kcG3I8+b3it7YqnJeMDUZDOA6vuhaWYTjtAGkSXfTGYoJHAP23JqeTBtZU2pZ34OWb9WYB3pL
5ojCoSOo8YySFPXC7dB/S04xvjxXJTP+cfPIG1huJR0YtRjYzBuWabUhsb6QkqTXDe3Ua3k9QWzq
/wfALkxoORX9H1DbUM/5q7n/rhLNojzMXLUhMe3X3/zvG5oI14eue38iBygP7vXGrZbLwK1Iuna6
8lrQyYn2h8+3DXiquMxuE/xnpKm3f6C1kicNV4mMdfrNmtiHvg2dgJPHNpLdqkMhDmLATWPeel1y
VEeAU91xWC/zl8/ddjC/3L3SHeWH3fn5+sSvjdooeumdQ97fIw6Nl09VvT5hPggNxLq/mNo29ti5
NF9KdnEKI2twJ/9AzEOkjmcfoSGUbOtZzTSVHGVFdzXD0iYHv/iWbycL4m3CoRTwtFFL1RcjoX//
/4ya9LE9iMHJifHW1IFFV44jqYYE74WOU3p3BpUEEFIcoYhVWLhRnlggHViu6eHvu8KLoN1uaBrX
3a7z36R7xus4CXVraCoPy7ZyixlahGq92p3kd1kulqkt34I1I0uoBoVeHxBBffV0uC++wIvl0zNB
Xxo0UfNb+PemVrRoHxwHvnTsMXxA/EH9MuBU7VsmLnUIQHlCqHqt7kALTZ+BjF3/n5T8escIbqNc
djq5o8BMCg/zX5oDa2CqECVnOv2TrmAC9Rd2PssiwTE90Jak+XgK52oj83HjxeiOJOUXtj5Tm9/x
+2uJ4WOI8FKuQHNOZsBp/mE0sKYEfin7ULWRbdlvTUz8TuPgmLiSoIm1m7ReH4Qj7+90n1aPG83N
5J16aKermpo0+4aFQ55n3O66VdxfsA1VbbHXHQHf4FCjGvca1DAbvaoLSb2Wgzrf/gk/afTdEYxg
k7aFMBisQ1g0UEPoRrxZciwokZLQyBl78syJAi9rO+/l08ypsQIPOj4Qzp/Nq0J7FVyBAwS5OWQZ
4muIjOx0sX8xoakeW1OF3u0gTXPRSK++i44cF2aHrkRyO7G6moFCxGlWJoALYHB1b5N1H2KY2tm1
SFs9XqvJRGTjpM7w/JjEwcQ3VencOQ2yArM2x+NYIPFyrzklcJVhJgW6FZNJpVFLi+Ao3mLYAzZl
pGhHvbwHpyKQGqx0+AJD3Bx81EPc7czuDCooVetHzb2ghVll7CMLYKloPP7BPwe9J/iUWSaUlz1R
LsQVAmKzCVRgr7oXtFPo8wfg6Yo7Cr6KCo3DcvvQNkrjA8k1p3dnCnsfmwU+VCj4esdy/iD1ebPq
YrBBX3Ewf2xOArJWFJWir2A/AFRuql63vy1WZXj8zOJhx+50w0TYEl0i2Aoy9POh9GmeYZjqopLc
loGOuinN98OhAruwz2kbzZSAzzsE4IWlD/lF6SvVU1Mcx68qMY+OeUNNwMIL4R2M91L4+nBuEnVD
+s9yFBW/ITh+ZexIzw7IfnaBOtpd2PCameXhfcOUtJfWj3Zp8TAyQDA1CVrk97uzGCUo7tUmYokQ
h0KoR3vNdDum/3O7Rv1J1vqJs1fbcADvgId7ivMByd+gFsWcfShM0/s78muJyShrSA3QZ3Pd8iTc
w0T4hOdDenl+ZRwPBmFIkBXuoVlt/2zdd35hBGmlcYayzklhrEGc8YHbvUPAXQxmaPzb/aOH1B/D
IM/MvjCfi6u4ybSBVz2HGMIMn4Gk9csjE8qzPwh3QKa3GjET+IdC2PvXnYBOAXfENk/3F/cdG16C
x/NagD4sytZ2LPNFXYhTEh3QaYhV5KX9LHA14/JHYBpDXFiO8F8gyB3Bnnsjn+L0aguP1uZCTtd5
jUFfGobhlLJ0qayn3CC70X19EeqT8WWixN0i1dcT8jS7MO725/OTDfoCPakDeuNrfn9YKKpZwh44
cIZ0R9wjg0A/Grwv/yOn+XJH5xquUh0F878m0dhKCF+UXcdHQpnx22LrndkAygWBZs7M/CXOb/aC
RYmhmK8y1s8GM0chkF3jmB7f9oLtIbICHep+Y7Toy0thPNVWV0P3UX2zaoZxbD6IKWWPDt84eIFy
Mqd70RTjFuYC+49mPz6w/CoJkoi3h1zSm5fKVf3GcrSja7Z9e9v/E6fPyAv2c8puxuhHOiJZZPI2
vcct+vsIWaV/mEvB0dhRIQMKmd1O9QsdRzDddkOBnPmBnNdxa4muCgah2NqxrOqXa8KDIMdDLP50
YTODbGTL1DKtvigybcSMR3zQlIMcUO3+Ye/ANv00hLh2GqudhPJXDDb22LHEakGRCY1JRS5C1b3R
fJmn3D4A9ZDFWBC6vjJFLz32gfEq7iNZD3mDW7RgzNgPSURR8+Awp0VFMf8i08ntutn6vQn/V4nm
JGoWO1d2TWHUQYfw/rzA0ERX+SDnEFAopCxOXMtSreWuL8+0UUrZhnsMSWQ4MAtiTKa9G0QNGMLz
H+w+PlDHdwwEzOtJ3U2YVyJr/cJOnO3+2P7hhgF1GmifiaaTV+Mrk+fXITR/Cx10ubToUfLMU5YR
9/XkRG7p9sANnF9/EdZNsTBTOwnrk6hNNdtE5sSwyu1LK2qa9c8usPrIkhyHBbRykZyEX4yt+0my
J9nPoygf9RXscyhMYrhTgFokISejEovPuDVRZIb8EYZbqcE2e6g+ixgKRUEm7gq3eM4SpWm5UsNj
jzS3bMvl8UfR5UWsg4CYwextt5OtLuUgDwZoxrdBru8LZVDVXakrLla7/b/fa8iNVqCar34Wv3mz
DuYsZVnqTiGEXzjTxJBb/iLAqwYRG5WdZx7weg6/CwENUQEedN0v4jNQw2iOaXrF23D3ir7l4Arg
TytWclzIo7twE2haWCSJ8K/Y4xDkgCXVM49AddaMWGb4zWPBik3P+bUE5yJtkLFDyru0ZNkBYrOu
1x9HVhsDGjS7cNgwgSDPInuna5RAUt8A3sRGfMGcwvnsNAzYUIGXxDQDoG+9/+p3gh7jcS/ys8G3
Uas5HYJznLF9olVz29ryrfgKAYNC2r57ilsmM/Svb7TeQg7OifzPPSDCf9S8rxE/ryYJqZ/IhAz3
5txML8h33uhJnOoX6+FrEvKjUogREWGJpRKvJ4teplrCJV977PTyDjQkk7pkyFYZCryFdwOi9zHm
OtaN5NLBb3a1DUlpIzO1yG5xOA7tN2F1+aXNUJ6PMgQumRAVdc1gzZrs5sPSTQaPocZ6yHEbQ9eP
AqgbZMFslgzwUgZiYKMJz+NsYO8gd4KbMCgB50/k5iKJda1XAMkpktIIlkfcbYOgvJ6JEg==
`protect end_protected
