`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
anprbIjnuIHISvJF9xhIpyTU434rZQIyY2T7w0qBu1FONcj0qxv8JENCWOTPao3avP8JQ1q5vylC
mEdeZ/EG4A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mTtjyYnsIgiG8BnaS64lZwqfKm27U2+ehY1w1QU1TIFrzG2utR/aHJF2rTNpPer1ErENgxU0R6Mf
xhfEs/B6+SDFTKsYNFc9OuNFcoPO+AoJ/u14o/7w94fViqlIujQdf4uhJblcVaxAbC4zn9BuUbnn
GIjAVCpriijhvoXcGtA=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kMcwwHVrWUAmpHB1hZpQeFGL6IjSMFRsgM2wDpA9puCtIDbpB124SM8XSjCc4ISkPwi/q1n3DUtI
3ETjZ+HaResnf2JctlK7ypZ5iiUulZoYRZKu7ubcE7GJu1ahRaSjNU3UzSErmeqjq11/Lb5nwMul
7WW0psCEH5R1qyur18I=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IAbHNgay/GIWCDSyIwjkLkblwmHaElcvj/8LIsKN3QlsrIXRl0Uv2qUujaxWmhW3+qqHPxx4kIeT
p2uKX7CMP+ORhnlU8DOYUjRveYgVEqPP9GGcLOJI5VWBnnMfQ6Cj5bqLnab/WAkBrAA5LaZHgicS
qOmV9oP0LdZ+U1KOAD5/oaKm4GJg2AzO6D2R0cGvLOivImfaKJ2qCast9n4RF93Kv6IZY54435P9
Iws+xXLPS64Cvfs+tvZENs3dGFB8R/9+lbe+Kpi64O0fVAC3MvA3xkmr4/1m92qP48zzneCMDyB9
prjDVeqa7KqWaVLTOLcgEp01nzk4otvFjrW8FQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TkM9QxHaMk7oZ7fmjKuHhIsx6aah3bQeK/SlmmWQXua7DrtBRuI6aWwWC3wywM3QtLCu15IkMOre
f0fsVilApJXXbv0eoEwzPM2ho1gD/vUWhitPHQ/goIBvSe3J75o0Sxr8OLeEfstIBP+/vD3XS8LA
kOKcte7S1g3XImF3TAMCnKUDk+OPGNVsJg9Dtfy9QfdtNG+ZdcuNPmB/d/CxQ1uW/eDx9gvdMZbg
Y8DQQ6xiqf6Uiy/I0K1m00LYU2/cxqy4pMeqi0r9OSOW619PHsGQs7xYs4/VK9zga5w6tpZNq2Q0
kvJWaTbdqw5S6bw1mu2k8F2la0hGRimITQpDOQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TrmmHEVLCM39ek/cnDXVNuJnElQOMHF7eZzv+Sn4fqZoZqQRSSMBv3Bkn2TMrtm0af3RYw0xKFzt
3Ze2HbCp+fAWccGk/WbntQoSj3cNS7iGEIl2aCcs3bNYQACOY7vJSjAH/nd17lIdzbP3IfysC7pz
KT8PEJ4WlW9Y0KygDfCaibIVjJj5r+W0dRTf+q5tDt5OPX5C6rkJhZEAXyJLQ8N0g8/SZz2jHher
MxgHDeB4BMeKZWtfMok5dUMjODIKJPmRqBp32hYHe56yd44rZ9UcrxG1w8zoF0cquHWujXR/Mc9w
y17Y+8uRpzYlZ8T+ujwXf4UQ87ZfVUCa8KgIzA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 637968)
`protect data_block
rYq6kq8GcWFlo6R34A0ZfM5UoajqxqDfflE0wFxsZP3VjJq1PkSpLXKINlnG4d6Le9Qft3UqnLnY
4YzfrfXNNYe5v2mcV6L2SATAxX33YOq14bJXTYMmi6xkrbBZKkTp3b3m4uTJH/Ohc5ki9+uk4GUv
AxAchipOjEGtd7yxNf/wirlzizFGjbqxytC+9pS9LdMuvRSnMeu7NUrlg4pqi+gDbFPaFr3bWHJt
J9VBuRUUIYqKc96MYPXn/oKcpL9X2OyIo5ugXL/8T791X3PhrxPUwPr9uxid5URLKaP7W+Lg0LWb
ZMxwJx/RusGyDi7D1a3rKDB+iwFIUImJMBwi8fw7xNlf1jEqJbcmDacw/+vj5OL49fTmYyNkC/bh
fvZrPx1g7KQVAIbkruHBaslVEaJtGYsqcA/14R9xYSxzMG6+Bk0Oz8AF01xqVG/rQbLpMKqA8HCv
A35ipnnhG5AW61foEMAG0CICkeJIBSvoHm5dPFDVYBYU8LyJDDJYibU4V4smQXpI1xrJ385THMm+
FDuBDaFqRs+J4/KkslFl/LBlXI0tcpYbDOCDxmPr22WBvSscjPVU4Eb2Q9pE7Fbsf+mlSIL6Pwrq
wiF1q9PaWFQTaqRU/MVU9J9lCxAVfzt+N5HCa8CZCB49e+ugwi97tJ7ms+cK+GqWiKbqnzbNYoDw
S3XMB15i4dgXv/sXKkSShxjGx7teJWcvXtmJfJ/t4P4TnS96fXIua1mT9tSTbPLgzhJAT6lEo2fs
0tT6aOr7nQkuC2/89G9xs2L01G4yMIuUyMUXJ2k7u5LzS4iiVeryGTOKPoX66EivDIpYsnym+s/i
6jbYm5BJpmVJjn0Ag6+MBLB47aPD+mredwwpNo8pK/B+R/Kgvn2vynJrWuZk7pw4qqX9W82Kb+f0
iSqYe2T6sdBQo0mFlRZJU+xCTAaEl11wB934r5b45L+4uzZIzzaHEDZ4pcsRSz+fTxoJ04k/hY4P
SPxMVlKDlPv7kQgdHwNaUzNJ6RSFHmlYA7kggYhipFV5XVovzAYEBQsu+zN4bl0u7gDlxOwyz/2w
7ytx/nQR7PxG25klD1jOg+UWNvielIVW6adwVEPYnUJ3J07wkdpWtT62jw15oqluWIsidnJ9rGF7
DyPgukSz4WvFRx4Tq//SNozOKPYH57p+nHNdHx8QxwhAQoVLEG+9E+W7oFNW7aQoYwRqsVoMOQeV
Dxz1vIpNsfWUUeIgoK1hccSK336c/i2VQmyseXEp4m6d0xXlqIXY8mKl1SlewZjd6j3ExDU4BdGT
HCMBhSqbG/VrBPj/RVTd77NIV2mKhP4CUsUqjKyYnpDSaJ+ZIRt6wt368LltvAbGaympXr9jLp2m
QkWAdaky3lTiith2guVXEK6JDXu9gVUjiSaOUBaY9nOXBl7vzZB/2Ey0xVlcqLADAxsv97xSm//M
ezTRQOvxYWUjZ0J8cGq302G1d6wKUrkKhQuMVtaZ+NTlXEd0G5uQQQsz6FVNxhgfnA08Ywj+ThQe
IRQK9lEEZ4U7MnT0nicMOMj1r7SsHUwLA5kLWgc8m/NV8yDwkKIP9JBM9igQ+/a3hY4vk+iBEgkm
uQLfR1KUdtmT8FVFc30Qi7/D5vrC0kmJa9Uw2W2qWkk9hINLpeZNa00O0J6lo0wpGJvpcNRHpIj/
mZ+Lba5d5iL0+iez38AZ0dtzRiNcm27BxqzQVwPksldBRB2q8LBW6Sk9Ua5GQdmjaBYECH3qEqiy
5f7zobhX54FBUxOU8zcTA6W+pJtF9pF7qKL1v8/+/I1/jB1zwpKONN5GeE5EpwFApaI5t/C52Fv1
dSk/ZAqsvTLmc5GPKRt40iFIKW5VcjfOQbjmLmyzhD48ZW8XOg3WK8AJgM5f3M9KAnJP8xbHULPY
7Slaqceq6EFE1TQq0SWO2esTDEaCBUil1/cwviGxKwmsGIx7Em0Rdj0bL9wbXYZ9i63KL1PLDN+g
bDvzH4zpfP0E488zkuGjz/SDnrf7Adc4QCRZ8dsVG9kdDymsAZyd4bcNmGWnLT14DzgzP9NjWlFg
5XIOL0SBfIXakBulJ6Wo3+kWguWSzYJoGWtUMw8yC3ai1221bgvoykDoKlTlwGRPtkNfQz2+fHsw
phO1SqxZT3KU/mF1za+LJIY4Efx81BK1rGV2LJpoPvg+pc62lJYypaPVdkWpGxXA0Y2qLZn0pLz6
qyr/4Mk9WAgD+yHMqDPod6Dq64B0zBktdSqep/US5bJGKYyZ2ecDXk2+INTVxZnpW3sEUWhT1kxq
SFqx60eRUAityYMz/XzLiQjBCnvTF/SBhuKP2Axd/mXxx4yxxqNZW9zpGc5HoBcUZxH2dPgURc8o
wCY4mH26SntnZFDBfw5uaZKABOElps91O/A//c37PIWnNCsR6AuDkJTQB+wgvN5j8CDsW/Ytiz6M
GDlql9Zgllra1bdkgiuhsna8u6a7NhR2+wErW6BpaKIBTpYOskpaJ7JlaJxReAbF9Wrda4N1lci8
a7KsYXHOgo+zB8Z8bvKKhA549Prr/P9jxTF13mQInda7Bb1dDj/UnDaakBWf6maSIQnZzSltrPn7
YHyuA/75LEm6645FAZdcwIDvtEilqMFYr82nnaz6tv/HQuEDDqNsAX0mjIW9eFAtunCA8tF+WQDn
i3Z1UuvOTWVkdGtTTQGHePa/SQz+GStteNKuzs5HMDYehyXQUHU4XzH+pA4T+NCuN1iQR1xFZPvU
8fcSioMEUmJpgD5Kd9TR53eEzM3TnRP4IoLWLfyDrhaiZzyBoWjF5mtIIBAqWCfISX8CAQO+JCZZ
sXoZPrEMeOsuq3Yk5zDvzRejoNgOYy3Tzoy8ads5K0fcbP0dKUYLIZwUgdU6LWzrsuVn4ID2x4/S
wcyfS0ln07U9OSELIFwa9JqsZHwqjtEkVXD9SSHCUDMf7vvfXwcahVzBPOsx/jR9eBG2+GIUF3ai
MrgUajZrfcTg1OSs/g/Rmxc33mmN5E2RdoxEtnDzF61k8N8+31aww9KvLRUTPpNtYgOcd0EZJO+B
VJR1+aaNYDgAYr+B45Lj4VW/rsXOP7Sb3Dxpz+TyYvZ5JTh4aEBV4e5PG1QfnAgzebZ4hFQK8P7k
rBHui/2SDbrJ9c1uuviWdycZhSGMV1RGw3vQ6VMcYi8rWlFjlwkgpD0g/DRjtgxRiWJPiSojjCnV
sCJNnNNKHZC5qyGld36K/w/X32wRH0lVIGyyApvU/yIuYQBRwv/+2HJ2Uxxf8TcFIKyasBk95w/g
syr1POWg6XgA7U+DBm/jhLHRlQWj7ChThKiRPcZ6Y6TFV2XLAAJL9TKpIKfZIksO919HJPGJGADc
uyWBG0bUzmWV2AGE0406/n3evjxuUcffuKHprQpblYVgNGCNdbL0kDnItHhaBP1TvGA1pRtKqEMH
OV2qXcbWdeT6sSv3K+QLrDH1v3meN8QGqhlboCkd+xXQXBEq4HV21L0RNAqz42jgwp0SYa5MT1dB
rPBo4IGwsskmtIClZ3aHC4RgmWa25UK9gk40b/72nkkcL29LJcWf6qWKVKDrfrJfvRjTHqksTClu
3KTghZA4kcsrr5/F2koApCDLu9jPdVuM8pyeon3F5Rdf/QgBP+Vh3K+0PUgNT1uKeN4K36kFc5W3
mj2pCJE3LM8qzrlSngmOsTDx6GjtwuPT+/eRWsDroLYUGta/o7p3pj6PZsINpIj9N6+Fems0U2rv
y7eqqwL65Pw1rolrdmHld50OK25MOk61+kyagIfTAAkvGtM+4WaX3SxNWUWct/uJdOcdJWzRc9bG
b9j4N9rNLTlA9oplCcXHKtWK/GznJrZxRJDdcFt0cOG7TLv/DGlzjE/fxmeBiICAuBy4F4UYYc/Y
1FZGB7OzGkcMV654+MQWx/ulRljljNdofrZgUtGnPQpxhx4A8WJsKtsOasF82TkSdLmlfYDdzqYO
bwj2EVrZsgeFsJmKVUGz2H1VWz7beuqdgd0RhfqFdrMnu93nuOH+R2ZCSKsj1vfBmJLrFIS2DCb2
7MVzCwrhRiFbQ0hNFzluVCfpj8KytxfEtEZXVcIZzAe6WKeOa6hkmqlaJtHkkCuBdwAYsTsx3vef
0oDJgTgxLC4O6okBkuDb0l1oXV6zzUhfyqJjFuZuheGfp30sLNouxfftHwOjzFn5PtPU/H85ySbs
RBNnkERZM2RetKtmZqiPP1dfa309flQbiV+CbBuU8TD/l7/a6mSf+iFhm++mN142H90vRcfn0b/1
5QawZCQAFGGO7tPPRar9UGGzdYO3iRws1tY+2WoszwNaY3RqKpBV9Pb8KoCXjZEgYbXuPm95gPDI
xrBa3zux6UirMmxPo++Lx6zEod1kF41wrs0yyk4hA4B/KM6l8QMIBHM58HM9o4brdpctxEesEBqB
bBCf48mFyacPtR1uTtdrTrZO7SWs3RtKDA3cIurWJtyeR0KnS4PDJKP5RAFQly95E4MmpEiKLxTj
qX4R+KgClCu3Gfz/Li+jhjbkbgixRAJgdGLXtPIxASPLELIFMuCqmrNrBuKED79VKq646YLYVF/K
hP7dh5GvDAW5KHRqzlF3OAYvdZ20kBhC70p3zU5igWBFTmuojiZF2CB0+yUbu7W/Jwc+RO/oMCJY
3sVSRtULEcAYzNPZipPCiKVA6w1ynr618vhATUlxE91i+YJ2uZp0FhG+t7QuH0VeuptFP9FQHjhM
8nUFA+9Ec/ZX+NQSDbbdhlLuKeN9oHkXBMChGQY6r4XEoGo30bRAyL5tM1xh7WDnt7NXx2b9DXwh
lqCDfsXPVrqGMl9orDf4F3p9O+rQujO6vN89JrKj3EHdmf0zzi2lTLR10Bk8wj8EB/UFNFHZFLKb
qwXyYyc8NmY1nPmG4jerBgMxaBpgfLR0yr5Xlf1rzW/UyyWEPwj8TFqsaS9BSwEQcMUt5Weke0k1
XGGHGr1TG8n1OmbNlNLwFZJHTS3/+vybqT0yjZTTFmv7Qhvp55doFyZ1BdDccQUY6P+Hwc5HZvLm
ScxyH/5/RVvk0cLG0xbcrekxEKaqqSxSjE9oaVOjUvSq4HE10ILPmHyzVpyzhB77WySnxuxr0/Po
3T1sXiiRzFF0MDxR5Dtq1bDsAdSnLCKUauDRmyXB47d3PXEyAD3R0cbMrM4uVylQ3TsqcsMJtuSg
V+1aMMC/AdG5rfM7oWehO8ERiJf6gqBzu3Mg/GW7wmeHF8ID/xKGhm6+famARcPbWH/phB/o/bYQ
JVkQOIwrZUtqfmMKs/09E9EVtyQ+AQ6oCHxBqAIZGHhrKbYdd3y7OoEJFt8D7CvyyqieUy8aMOPd
DmV4Rx9YIVoAgcJZLFqB/+eToCAfzFqNcB4POrPm+KIEKX7WRns6KwQuuNrIBtpCvt6QFmE4BU33
HL2niPXPikYaoeqNuhR9zovrfkojFzB+d/Tlt8fwS2LtqSaCgmNc8nZ4Jz40TIC8BASbPcwN1WGo
cFseAQ+ILq6tkbaTsCVLYKN6B2z9SFyr4IIXs4HCAHCk8Numc54/0zKmoOpJb/Pc0xQIu9agzkMG
C4QnAp7B5cvOZ4KDuzXgzoHyG2pMXjaFZnAoaYYgfYpYeyRRjw4d06xNy43d9FtP0ONFRJvXQkaH
4IApa0nM9aUXOFh1ieWMHwFt+saP0+EffCcgr8fpdCBgBqFPPq4PZp9L9XNRztMJL9gOCZNlYQel
ObSUI8EZp1uabvZq0z5zWHUd1zsQ1xg7m2jS8FhZW1ojy0itYB/566ZeZYuevm67OBFfi7BXFbxc
si7eIPgqGVV6C9FX6B4lOP++PhtKcPwVaVf+WEisgS3upWvaGuCOtrjsY+R01cz81wLjLyOfRoSn
+Wh/dbQBXA+La4Hs8qWFqEj3tq+/+XvnlCjhmTyFahKi5JH5oWS9SgLiGWX5GwJHbdlxeHhzkIEv
a9lp7MschR/iw6fl0Psv4loBqvnb8llAnVHis6/x8LAozQcRlKUy1pw2zv4P2W9kcl0lReQhq4V1
JMuh5/j7EOcDpEojQBtYXVdEXYSDGhoIX8ljA8W7J50I/thoIw4F8HiDYzJ16csVBu2c9APQ7DRJ
f2IZHo4jVEjmJhLWNCq8LQtUjRfIpuoGh/2vnHweJZxvht3XG/cU1KkHtBWxsRdnEyBqET25cSaM
9lS4HunF5e3CIcNG3y9LlNRzLArjxVWKo9I/UYqG72wt9drGB4EJYWiFrmz6gsbvRsBgKMD+feGF
XN4ReOon8wMd1NYgDKKTg46/jYGyqKKtquQNlZr+TD/+/BnPwf5BexUc/mUtHpLr3FbTd3bWSn5/
t6kuR7d7LTV0Lxl9ASrRiZN+DUH3sYI5Y+egbVAg95sUGSnYAnKffI7EJDgI5o+iDQAryEW/PfPh
ZKVUDZOFRcOfCGFQ9S3PT17vtv72jSi3IdGB2heAAKIO+iOw/rax1kueRX6nyrI4Yn06jJpwA29U
ewOXwByuUObTyCNHD45tSi7gpulaPK7yn9XbpWV2fyDialQBOHRihD9hGtWk+iSEwhOvjTA9sv+q
Q2U18HLTGXd+udPQgkY8ixQj1F5tOVcS4N3U/UFPBNqgq49DDVYstLvdqkTp0ZA0JOTR+ow83cTX
5LxlM8M4sR3y851gDSkdEoPz+JADF/Th9TNa/yhAVy7+Ea3/yggAeB4GjlzepuNgAhbA7QFz7Qt5
ycJV+TBpYuKTJOKSvMrogrFELKQ74Xe5OTaRzaGXBHI3+ee9UTBF2mtGhjd+DVVWbEanD9I9OZTe
NXhQFKh2B+dGtHseq3U8lwlr0SQ3K5XEuRvyYc6LcesqX6W1QFxoFai4y2KJMAv3CPs3P8nm89au
RHFjq5lYID1cmXhuwjz/7sniGod7Kgsg1Jwn9+VyX6dmSShUMtos1WINmoIoB/FqNZJmB4E5V93b
P539qXAzHEUVJnnMNvckqSxZz4aHZ4XSUOoQMBiS0dKC5w6fYlt4ljcdyNgTLc6B/xHmK+hMBIt9
k79K1afIe4vHN37xXOubxHEnCcXFnfm4ROGGOaISahaXd8mShVjJkwrV3X4nkBWEcpqvsVJ5+Qu5
herHN8pAi4Gql6Um4EC41iVxZjTSOLBauAmhjaWTq/mgqmof9TSYAtBIpJq80j2JprMCeDsE3g9t
VLWwKmlai92z3v3Lit92mpDxOa98pZv227sIckC1dLQGdPiA5VlaCY+qLI1DzV3+IZ35e04Kz8MJ
/544bnPlj5P5aa1RHSl4S02PAW4/xAOT6NNUjiHvdRADfc8nqpcWM4Viq/b9oexpjiMXQ7GXcieX
2FLrNvumLj0/V1i7wGXzvreChP1PqGsnVeHhm2/3+iIFMez41g4MhKd67IOq28qAChUvj0B8BPEn
FclQ6gdPVOXMdT+fv9TWNHPPSWwBkWdjR5A+XSGTwwYKs8eqdURqDFSezzXLsmuVNJi64ScIY3Xx
yY/p/MJIuhCG7iqHoKLbNdGIh8vXf5ssEyTpnvWILptKqqg6r25Oz9t6mVLdlG7YGdC3T5ukLKKv
YP16l+l0ZUzYLpdUcU3sCZZumBS/R1I1hv00cZ9F1vR2HYJ8SUVV7rjEyaQK8ry8N+BXf2WIVE7f
0VtBDnaVpfTPfnw8Sp8pt0LDHQfwWtfcPNOUnF3u01YXb7tzQdkkQfZWtzlqJNtsMTj2Tcfd7Idr
Et4a2y2DJ8o/pwkh2D8Jwch8PlivusmUG03qS5x0jm1G4mzeOvvfkV379DTes0KJMamVp4Y6sn3W
fEsSomcXd8PDOMb+XphFkB93gYg/IybvRuBH0IIs+1MMJRvwdU2dOU9757Nh+8AWAK9Duz1l48No
oi/l6D4FlmvhXoU26LRA/WpuZHcVsEn/d8tS9GrulZSqTZ6S/x+W5NxbXM1soIQbiI009JTVz4S1
P8rQPSkDQzLWHI4+IUae7o2vP3+cMeUJVUyspoByIE6MitZHnheq0TNY1L1Xlej0HOefuuqI5Si2
mvj0xntCdShWwzPuQ96L78HYTHdwkVp4l3AGLbOXORYWmH/IJgA4pJpH8tiFktn+uQbvGTlQ1vEG
Z3+j0IOn4/vxwSFfwk6ZgFmjGkiZBdxYNqroL66WzaxjuXE1Pgh2t7ssVPAiI9LJG1Y00BTOz2+w
7knxfgvJ3NKCSZOkZ6J0Hsx41UipJkjKUWGDyQDRg25FmDtlm7nnZWIRKiS2GvQXJoQBeioDXDpH
06xf62781885kvl1+EA/axBpN0K8zTehV7Qns2UM+SCKFXJfOk/ttaBsjJQ3O6rQxJU6kYLatBPE
4+X6DoaP2s+apmSlk7cafCuillKPTbS8lzCPuXDjwwkSwMI1CVtwjIxojtaHSQ4Z9YjvedArulXv
AUFRPQMTf5EvfcYmQTYj75ImKfNZQwS6mIEgmM20PnxuoBqgYoKEg8TCZZEiuC/lpDoMksi/kQ8P
ieVda01+1rRgy7PBgsdWWZU5DJyIo2ts+RnvUfrFqe3AMc7YA1yoDcqR5sdy3KTdeHWBljQBjTg/
Ol2tTHSnSUtPif989/m1+VlXAc7ywTEB/JjXhf5aIyXtN1nctYXDZU9/w3k4lLIfzZ0JwWqPejjC
72HnOSdrsAbkJY9cem1qZbsbcviIR3PclWBrRcfiawoYYtNyTfDnCGdzRRONgWP9Y/jUaVJO/jk8
ClHes70O3D5Xc3NIcZErn5JC0JqtSAlooi16Qz8SmIH5v1Cx6eeFQi6EGLC+CouDWM+/1bk41O1V
qfvqDf94DGuyj6dzKRnyHWKGyxOMyml2XOfVPosogWuFLTs6DZWTpunaSRazNLNh/qVt75KTUxix
zIwCBo+qoeGGnvwHDEiarm2jUY0ukEJ/VHL4D8W4yoiQ0EH98hDUO5sWE5SplVBJKM96/g/ndbuB
EZPlmals/PzgVWjfhy+Uvqyj7X0PeFv18CNMxnVs8QxNon3cQzBzeCa8iUfzHv057ncEzYZF8NsS
oIcknQzTe2DZxlWvHc3oy2eBX/iQua80wO2/QvTn74JOnFFxFIGU3sKng6GEeNOHcIB1lHPjsZq7
5FiQWigSc5miqmwNCR7myFD+cchsPv6O7CFIGyk3hV2HwepPyvEaesK9ZT1QTwCJWCUT6osm0cRX
b+eDMZ9Bjps5JwR86r7a4X1VDKVe87JQ3X/kTuJ7LgkQlrQ8rY/NoyQjOeImvGfw1Ymc3/zJrn6w
NpVG8vza/2Jj6x1mflw1iiz98MTcuX2GRErgnlSbiMWORTJcYpaC+SdSWJgt02QT/UXx2Ot/HPL+
vnRoHC8Efl056SVslkMaXx1H51wNiMEarR47P61RS6vAkqY/a02ShQ/K3agk4+MwoF6cHMbhGg5i
bDkvQORx3UAo5epV0H2pszfJlz+I0FpHnbpAur0LypKopptm9czUZFhLwecqPG19sNJIeykY4YNe
iU5TBTyJvwGgttobkexPfhbM7Z4ZzTRPsUIL/fV62yP0R/LpwU0MxLnwRSIooAbEiV8lf8k6TnYK
1BipQB2dS9GnCEVTk42LEl4iAyxubW7CQphCf3GUceM7Ubf+hrIlMP+HVTrNLpQX/z7MNB0X/2Vr
tPRoc3fw8ATCiXpCfyvCMn+/XY1zR2TL91+oqlrtO6iVingIk/f5jGCaqWVkxWbSvgPn03kLefMB
cnYncniV3gqEY3euJtuuci0rytOZmYoRH7LD6f/GX4iCZFrnlGx52pE9j+Y05NJoIfEW3a4a8rGJ
r92RyaeU6yoLfWQbHeWBN1woFIZAcLO/hrm64clpakEt97ka4GMg3nRE4D9iic16qgSY4JWWn9od
alEoTHhP60Z7e4K+wmQ8vNjXUi7akQV/aW+q1OK7dTWi3VLF7pZL6OFMu0U6iN1yKgP9fkGpqDDS
GD0CN3a7Hw4vFIGtP1BZbfN7oZU91FewrRGZOTwFOboRlgEx1CIjxesZVnO5b/uNynD5sxKJvXn6
H+ROZJHupPqCO+dLt6p8YeHXFdPuB8xCYCaYri4PIHfu+6UPONPKM6n/VbaEhDvHXmXMAR6fLSvi
lLEhcCHBy2ooqJtPk+Z3JrepGsQjk7vtb8qAX3LB7/zvl6+pMB7DP/bNSbLGSeiwXcJhygZrMzV3
oQIEpTrIdwGzIJZ1ilFUJxAfxJLFrm5rG7WPVrnOH5EhCPU6SQPsSCqIsSIvOdxbO3eDxEdhdLYi
Ve8vneVHlQ90sZian+FyU1paMqeLo2X7mdBtt2A5lrB4ybibM3TCZfc3CVZJHI9yFvfhBhcqpuwy
nA6mhf1ao7zuo0Yc5q4mX15A/NNkldlUD/olZC2CYGpwc0ro4sHklhM431sCvrRm7WaSJuhmncKN
pUwxTTebj/D1yxzTKsYGaHYmXziqPll7fuTlkeqQsWfPFqVU5MUS4H3N5Hw8DgXcqQFBT5r1mSuV
eo7MyvQtz7BM+D4PYNyLuBlmqvmfkWB8dIa2Jjmdp077jbgtNCRfujfOIeUa/M4IdlbVowKWH5ta
QOevwUSq9iOa6NOYLffhz8gm7oaUDhcN+Xg9A5YVNJg6E1AP2IfFoLud2BTQpRs2wGhGW0lrSEUa
TLACva/1fKJHSXLoitSrQPFDm59jhwN4LWl/INXj6Jtrg2vYszrjxiQ0EQUJ8SGMLW5lT8sRo59E
XMBzJH12tF8YoBvo8NgbXL9n20lRQfe40bpkue55BVvjggD9XT5rOD50QKOorR6UDTveNsoOXxDi
fX3ZeyW2yF1M+vYBOYR/+HrJ2m7D/fS49r8X3CzNyIND6pgSDJJi34+S5D0NGu2r2iwVhAvvCzzS
99m9GjlUk5oJmocvChGSmdrKfhpt5yuBG5esUREwRchuaZdJVWc24IuzmDg2JTegBf8T5IjkrKiV
9Zg3lLYCFm5tzdyuA2ZkZFQ4Y35WXgvlYFBNfZsb9O5xGj5/iLXqgWSP3K2VIYxWKtSUUyi4zqCe
MShLmYfpvHYRQ5oqM33lnEm9ZQYGuLgc47yXV0dffs5zBpfgx+c1Q7SG3EDjD0WVqPk0zzERbY+t
rQjWm17Kt14WmpPX4efWGrVoLkJtlhl98lENbF4PgIGjHgqyzZJwfFEom45JYk5G3RU729bhS6uy
oO6HJkhJ3hf9GLv/bekguXPa6HZ0JXB0oN0NqKnWh5r6agh013fHJ7h1cxZxi1Vo0SrAVl7FsNUy
P2N4rq+2ppcAQTobiYepVvTobUidrrzbplD3o8h+Jde+cV5MslEsCvl8gfCrAS3x9ojSc5wsAFqS
20emXexJeVERnY65bQQl9gSfe0lIdF5i0cgGOHX2OwcHGsYQ1+bpctF8aUaYikE4+ztNpZMI0zWS
eEUQPYtV5yypv7mppAr+8otKZ+mQrnNHcNy80kWjYY0lCnAMRxtSTYP8Z+Z+nchCVETaItFTUpNU
r6NJjmmABLhmdzcIMwKqljCic9F7nZxJ1wzSjy+nOerTFe+Rwnh1ZxdMAVoqltQuAzexMvRYhUSj
E6q2ZUS1DqF9iZFVDuZxUKCD8k9WxtIlr/Tfh8SDbVcBiCem2pKHvBoOzQv3+KEeLYTPR/4qVWyx
t6ZfoL9vICT3Qg6AmSNbe2VG0SyYquPEuMF9wZj/H6VYzZtx/yQzwJJp2qrhsy4vU0ONHghyC+rT
lzk/bWQlzL1JNxqsSKOmbtwFb8nDMIusoxwud6IcWCVTqcqXh4efjuThLzXWMJndC1Vffam6Xcc+
1Xr++RxFQbq6kxYflgsgBWpPJHOMvsCGlT6GUYDRA5qQu9jgjWTSAKYJw4b92EqKjOjC0f0mxJBp
HKK4AuTCoRAud0nGaWtax/CcBzRCXm8L4aC5yEYj1GK2Y7Zc/kswi/frzojbmAnRcp8STM1DAdd7
ZUsy6+nh4RrUUijt3EC5Lf5y2rMc4iDQoHBcrXKXOwSDOtTN3bYucMkh1gwT9vqjQ/KU0eZgHwQm
uewXMjCV7m34dIfg4U3xy4V8PzcFag9me4F/atc8BUEnV86UiLbPDtBfnGqh9AjwCCqIixz6FFuU
eG2HxNoCDzuf92pYGBqVHxAS0WtNQETm859vp/fcWWpQgLcNVyYbwb0/E69NzYpp20c7bL37ItHO
MJF6HdRnTllbiaf9IqAiREWxaSqICnDER7ltfZ2BSymt/LzSLU/o0qYF8XsM38lBscvWq49DGSNk
e2W8omUeTEfkT1QbvNz/s3Evt143DxAZWyyKXez2VMPw0AGCKbg72sjBSaJvxEC5Gg7F9KrCE7in
lSRkcPNgKGNdJaK9/eWIxwsc4uXfSu1T3aJ7HgyVyYdBIEJd4O3NPmSMzAPv7bQoiVj3vI8ly7jv
Mvv7mReSTc1We07xGMy3Dus1ooOThK3llkQ9SGOSZPFfCql2abL4b0tHcaPCoE/1r5+uFpQqHbCR
XRqoh/jCZrqg/jrP0yGW4q6qKtB4hcV0x1UStoyHky1uvMdJpyh8VDnuG5pBxguGuzU/5r9Gis1S
7WXW7WG03ntPg2N2fYjL8wlMO2lrhdl4BOJPecOH47DLr/nOhL+SSDUN1vTuB8U/DcTGkVXwbPqM
20K8eW8YwMXtktb3bDeMreIgneiPyJWToXmXh9SkLZv2PZ09aSv+0ItFX1RlK5SvUSXoEZpYaXGr
f1B3NjZh2VZqe73kRrn01gpQnWq/gZnz8AmgJGEWAt2bx1p0qU5rkw/psU0n6UwulR/oSyEVbtu2
LZW2rcDsrbG2C0/9g/ReYpH1dXC5Xe3qXYNYhqq4ahsDTxTSAqBpa8lYf5A711Gqu/Hpxx9gJyNE
qHPpDKri/CN0keSIvJtG5yzkSyRzY9XzgdeAr6G+TUqM9ndUXwdDKeyYGjpap7bwNLejHEy2C3OW
Ra9auoNdn7E6i4hn/KHuUgOaSjzUrZjuzATusUQ55XNzcbYIaAcGx3JyWab1ozkYWA0WFCG+neMX
VHZhilYrRpH79ZizShKZSRcnMfXaBtDdsvHT/LWcJDlV2pj1FG2c1JAfxs/2zaEuN7kB2hrxmnK5
TQ/Y9M910z5JP9lx7F9POUXtr0MigmhRjnN0+Mwqay0oDcnxuoX40fLFWKzos77B0u1UbYOJxBcW
qeBqSUEeZu6OP2xcFXn/UOoxJW22w9D/TysrmbF4qs4NEaafh+9NrCgp/3lTYxpOqwu8CvQ/ZZiw
37TzlyGA1lFTyIoJBOAOVTh2ws44pFbSi99ciO1DbNYcUMdZaYplkUYbDoBQYVibk6kzm48GJEH9
1G+Vr8V5YBEgnIloAjJl4dALcPvQPfj8TOlprOgb3fNTQV8UKUlpkxZBJj4XhOHygl0KZ/YIVloi
5MRR9q0+49tGgViAqaKp8GlS/2YPJwJq57jqUGCk99AJGekuS0dUIDeGzj1dSj3KRiWIWPwG9EC9
cupKtRdcniFpvvR34oxbWxWnLeXDWsTUJgOc4E1Ynjkkci4Z2VB20WWDmAZavbrWjgFDpLj2SSnu
HLFqQqbscSlLGRbq6wW3d2jnKskEVmUJBMlYm8iqa8k+ObblkEHhSaWlOxzGMz5XsXKkZcTVggnc
aQLcEwacau26WJsGAtTf7Y3NqlBMx0JYj9S9zlEifujjaRx9Wj9xLKPEllRMIErntxAFPagdYdg/
Hl0Q8wn6uTwvIjlKf0pDn3NevrrL873EsgvrvQrjI2VBnZjrLD8ZFJZWPGam8EPduKLDF7wFtAYK
DrRcxu7Lk+U0NuS2eNO8ykLNH0v/zCNB9hcyM8Wf8ITFfvsJMLEXUSUKsOnxSARdmzvCtf8e1gat
4Fb4lEDN8dkMkBPImp/ELp0TC+Si0yrzHYAKjG/6wf6yQv4AJP/LrRZRyVYApj137LurtS+Uve65
d2q8qNkNmNOFaGUkltDJBam7xko56rcy5Oz4HVq1qeVU0xiKTSIxTXx+pMHtTd96Bd+ReojSiYVo
bgqsURi/hNDZTFEhu8k66sfbUB1J+kUyUmVH+KGhOnUTulNiqbyQ9NiSPv63MXkfmYOoEuC9AAw7
Das0yaeqYYgLP2Q52ZdQ8X9+ivFOF9lExoc4epW00AOMbih1X1QyNnp12hgHqd+IsWkHVbXom+WR
VwvD86jWBNJr5/JL0COKTOH2Kj9XEJahK4B1kytWT9Z3ijVQ5JDMA37UIg1A0+rD+51SbghDlTl5
/BbGHZKm2ICH+Jx6Uix6LWWMsOKdxzrSVHcDbxo0ohxk9QEPi9eJR40dUhAiM3ZAV++UYSM8mxFG
A3RzhRI4876QeiYQmUNdbmfJWwjrsN+910E5N85RQFFhSfZfDl4zveV+yDHoeAQgK8tV7YSwn66F
1BeP4Zk1Zva+sgfNAhDuLcNuTwvbmJ58ZM6qRBLwyljBKdQJbFwkt+b+zxISgDmIL/2pGttNaXUm
LcT12GS78zNZj7a3F6lblNc8Vg9xsxcr8Z4lYByaw+YD3WolZyETs84uE1rA1fovYT9YL6VeSqp+
W0SRe9jqXBumUHk0beK4M1e3ADuX3J8Ie9pSchf8HVyJ3Puykair6UENFsxxj2utYJlQUNOqGq05
bWXYUalPfR+xUoR+KGvZXKTbiJYa1LmXCkz26VCLUumDHrby0PT2RaWGJzyLVJOT8qR82Hi3lpqh
8ItRhoQj2rvJD7AuS1rvEki82aChiTSqfrj6MquydRPHo5JCgtKxHCU9KYRSZJpcM/V6mqWwCFSr
32S+atiIiZxS0iIqpKOI1DytvbkxJaVlzzvlkRqElGrGBBnLnbax+nBiBhkcWA3N5eOeuVPcHtmL
hIKU7t2+kQbIFCse6mExlXmunw0A+wBi+rv1yhwH5xTCHnDnW7UuAHYIqvptTLX34g9Eqwj+YQ6L
vhuTG5ttuHIGhxD0LOURtWi75gQp7yHT0Gaf3XBisILvg7jc7mnV1qxdlHT/9D7tn6WGh1jWSABL
scZpaGFIu8evq62q82xNMG5G3DF/udWHfHmzObKtHd6sWHkZV/QbK7kPrPcX28CqULG57DAxqaax
HjBQFI9ILP0lHesAj4wklA3t2Sc3ExUHoF8Jvov8CSSWa8e8ki4/rfJwYrQ0oHjcCNjoTyR0xxIr
cVsk9Zi0mViagVIA8lBFnx4oxzTX4qms4LC9F40zXmbB7hQht9i+6OhSNrgYSEg6EvLHj7bvwWkU
q+tuqsN5qhlCsx2S43SUxzCb/jO3nT7fHNfwXFEgwCkojlobBiwbDKncEXQnFigLfy0QRLlwth93
rkh/zkdi709CEivzsRnxORnOMISF3OAYcZ1nAfCJiNA+w/Z1lU1YauEga7ojjsOFH7HDZZLt//dE
5xfo9eCzlXr4glbzsqY4WQsBDZAM8QNRL03gG4XrJ6reJ7WuqHNKzXVIfO/iqrEswIw8m4tr7QZO
FMzG4Lv8hNHo8OVaNL5ihvzT8vFaMFzfTNtxzLm2CxO1MjpSQ2crpbZm4LIvtKVkl3LJAzxVF1HB
W1TzC0ATmm1NRKRPiGb2QyTxEVEWnUmr4rvoEC/WB+6mHWNT0mWfoWLYLBi0Dvji0OSWiL7KkHO2
baMnWxlkOf28Ho+u8kK5zJNGX1VWyK3Nuc/8KmHg7GG3mgoa/53mElDFPatam1o/PZVYIE+gDbIE
ZHR7xrZQ1wXt7UpdZUFz2h5OKCXvlW5GHbCO8323bQuN2Jzvkordw1m6rR2qxyG8nneem9WvBPYe
1dxBjj6pP1A7knttqgZ5TaP8+cPp09AM6qcBQ8H5re2qSR03PYraI5Ez5OpI08Pl+Y967BG/0Xvw
1J6d7UpZPWPmNIz7eabBqnB5vo+aEyISfj+eMqhYFIdh60skDPP/Llx/uKUd9aysLa83qFwp+Cgo
qbrsMNbpTrNOb/SoyCp29I7zMtAkUNZue1DnktEXQ7uuDSZx13mOBYrxx+u0GFr+50i/By9Sz6Lg
AfxazLOo4sBcAzBIZFRzaGuXcYqXpKPm4gwKFaTj0uYd9NDwY3ZmJEJrWfiTQzPvIZAxpPbJ90Hv
RzzqCMFV9S1FJKzGXVeAE3+xIIL0y33UZQTazbqsUQMc54P/BRiJK+5V1Q+m5CKMJn2MemDRF2v/
uoYbdE2fhWe3YgvRXEMcbFFUt4rSFMxDrNtSE3eJGBxhzJeGCrqCQVkllzxvHhB4BFI0Xmc6DR2+
0L/V54oXgL4dIXT9l85wWSQsHsYZgDKZRvF8iLT+NakeJqIR1+61WMDwt3wJD8klRgznk7E9wru/
UmDNszx2vHf/MqdatLK9tY51P++P7of2a5/whL5VjdNEl7o/5wWTEaBo9fpJwLVcvr0mfHuaheRM
CUjCqK0arrtKJtY5rzAwD8pIv7oB6VJvM5swn8Kwmg/0Glkv4XNVvI2ozZwroS7lBF6fWNLv1Bf1
tTZzsJT6NzWL+5hac7hCa7elbaVnVibbxWl86y9OcqLwa+5gDPDPaekYESCVS+KQ2sSil6fFGbNd
qx0j015Gczy9gjK106hXF8W3b/e7ZjnvVXdUIfIPLpRWC7WcRvoLuOhPbYgIHZO9mYDnWWrdLnbS
iMo++Q6Vt4vWpLHwILgObUFQxg6wnVoKvV0zY4jMr/dbAhsbtRSowsCXCVmdPKkFXga3bA/BnjxZ
nuE9x1vK2cUuOd4Q/QS+EREBSCUUAbP8XvFG6LiORXRZol42U3iM9agaMwDEgMzIxbxz2n+9yAi2
5ucO7BVBBjnGBkECUmpxdEkgOqmWEKzNQ5JMIw+GUt0SwMbgF/0S9xVMlf2s/b/Hm8M8IGwtEQVO
4a2gpH0XMitcPRi4fSzoQHZfGUxk2J9++AZrbHyGwPjNUQp2s8pWi534tXNJV9bIupssB1mj9iho
g0HRrrkQ3CptL0v8+fzAl88NOJX9c6dmOQ6LZ61KAqlgpA/sR1zQLwOpEqjT3yxnTIvp646MXdB+
sDX7j4ligv/NNyjvagn89VDiogKGxc9WRk8YpEns4fW8IjHirukSgZupJh8E3Cq4Nn/dD402fSKH
gHFjj/F+3x7D9l0Kg2CZq1I+PRy4fzzQeQaBgCrV/bBDy6DaIQPDR3etubmwQuxooWa9SST/RcF+
u9q3JyJMtutS+9Z2C5H/zo0rbdKa+a2/RxoKC20TzyyAhLyQst0b8OwPGwU7aMK+V2VNoKufVfa6
e8FwUINxSNn9pxavXZlnc222x7daMJTz5hzOiEL42ayyxFQwJCAHPzyEr5t55kcpb9U0VoujOeGE
xGjLfZaZd4tZfkD08Mt3m82NCwq7QLLtFSiCaWhe9lslQ0HBnWI9rnWhVJUgABAZoNTryfG4EOPu
hN2Tg5F+rctsDrQwedSzHSq2UGLosiC0Ut+5rCiym1EylodL18/NIjNQwcM2+BcDExuPtbZkrhLl
KZXExiT+XhiNxYSRDauCQl1q6+YZv1PLrc9lzwM8XrKugJafGrHc1+Uj9QSlriCoGyAGHwP2LiJ2
LVjjcC5lMC8DlCVkFyFu3w7TbLYF5hAk3tmLMkZqywf6TuWkc/XeztfMAtJ5V1WVHndgmijAL4+Q
zm359AEYBuOAuzHmyiIN5RIOkvtC9h0gYaQ6UEMGRweqm3w35cTOSXXs4ReX8E4slRxlE9ennw8m
YO5nUs27/uNDA3sWR1snm92AL3KMzgvpbQ1n7pwSlSaLZb92aX+JYvnOxlse2Evj/WxBQKaxiwxd
HO0MqOvvnb36er80uBrkJEgzHLTAFBypStxqRh4fv6X7p2dcVRx3iaWschZbBIMamPdda6saDl0R
ESyFEaVzngJZQk5ZXcOZSrsutNoCpG2vUMT1nOmGHnUtaqV/VaHHJ4KbrX4eLpB027+yQ04rm2MA
AKlydFgcxmEI+qBPKDWiDM34TzT7ZNd7xuwU9VfnzMvXcNpKfMoNazRRBpluyWaRxAB7PI/AYsSo
jix8u9vWpas0uaGr6OnUMywNecFovXg5FfLWXo/S7UV40rD1+Sg39DBP72Rk+inxHkfX94ctgeUA
WWtbRpWY6juhyc3X+B90bwCbQvMHdObrKChIdgiqGQ1+hAk/uYusbybAcvemQijdCI9FKUYZO9ht
bWKcYIkg4r/XaHBxSCwuAba/ZXyFAAuLdl7EiLfX+tE38/2oYeXgSZMZ43DKseLDiQbpgvDqfQyU
VxCU7/twuIkAQdUhuoCYa2b33HJsm+2rzq/sxkp+YaJQIWz96+bjJoJV3Xp9KC+W0CVG2M0gpKKe
DmVM1/XLO63k92vaapzKfyjOuerSoTMC4jHOaETVbxLPA9bo02uxKFxkq56e2BqBkxtqXT/nD+Qd
KoS5aMDApORPRrgOw3BNWZTK1LUYsmBdd7eMeRcA7cnumVMnkU/xwYMwLb0ENEVPwfOBYj3AD6Wn
C/N7ybPAXwGOBBVzd8t7tejMg5R/C4tAkiCTBkuqX0cBrkus6yGpuURPxO7ou8JMnnaG863SqJWA
LASGKHh9C/K8W/rtTCkz9S+9MDP/9Ay3LgXMvved98BAU/xS8ihy9Xzk0re9Kj/jpsxZaSk6Ld5T
lhlcWa10nz9zUVFQoI6anlU0J3hfYp7BVw85XVVQB8XXlO7lv0fbm9TvU4ZutFQQHRnhSy9YiEPP
2DPlC3zVYZ92dBZ6WNMSVIB6mazEg+IMCyeCbikiY7hHiM6bAXgcAvcGZCNdNJEryzVBncPoEaGF
/fUxIMxHnBeGflgSkM34deUj6HRSctBBTfJ3Rd1Zy+Z0bi9hgM9vY8woeyHRm3m0ZRwbG7EOS7JH
Y7DIvXQSgjNEJYpYFb7b6vgkoCkLQLaBylF1+v+KhuI+Q2gsqcMtg1ZJqhaY14zzUIklF4ywn7TA
QdO0crsg+6zijB+yy+gZQGZSxJCe7U0XP706xNWWKcGlx3gUwa5Byq2RSikPNBqCsaOttNL13hj2
t5nJK8pFR2N+eMJIckFEFdV1v2Dq9Jp24jORUkIR4PX2I2Y02Pr/KIdm2iLpp+0gtIJQGOYx06XN
UHlroXg2u3aU0/XPtSclUmv1oy2d9Uu8vvz0tMMOm+8x1wjtNwd2fCjqy3FgGXytYPkmDcomxr+6
QuM4Kdd5RgfTee/l5JvnwQweKAMikhJh7gGsEE2hGfLfP8uM53RGzqQBfxV9Mr0LuNXLD4b6nHzR
Z1PxZrAj3teKHNrGRIi50SFSJj5AgVrpPdBFKSDYGdw+XtIqLRqSEoRC3C648asQ6rrN1al8uyGe
RF1E3rQAVrMbw5iWcZGqRBekWfPfz+t4g11lSy6lLyr+L9yMsgwfhMDLwo9s6YDt/FQkiCEcxFiZ
9ShJc483ooyA8e5vlj7OtiAUt1sPCFrVvqlT6o5EwYvcE9dCKefrufX16tsXT74W+iZ0nOPeeKhH
bFhqHP8GwtGbcMtoUgpzQVgSZpTURzDBpvM4iWWOOLIQv5PkvibldOQX1b1rHjwpilaWwEe567QB
nDkQJXjW9Zd6Hna1WtCAinRUC90Koqq1PO2t7TlI5Vjo91xE44AcgXSD/bxts2uN4J/seYq9We8D
r5F3BuqfecsW22FtqG5h/2NpVHLcVHPIOrBk9Ll55ELJknCNmefor5gtz043BQGq+u8RLm4m9Ilh
Rbi8ip4yJQEE3LAGMmHBo8T/30UIwPMIEkRbmvEpRxHk2dd8TBXUbo/AzPPeZ12RQbPNSLXhClhc
Hn6MKnxxVLTLJ970AXk5EtDFTWN4Nu7Wm1Ti/lP7rqf1ctJ+ZO3plvXXXAqX9m0StWKXExRsjUO0
hm7lsuScREGs8EndrlZcOoqmM4mTjwpiRjdKl+m484vG+glDJx0DS0OeiOJmXjatySoYLnX6CkjE
uRjnPK/stt+wEcASZrpnaDlSEt21mBnCrpEcPANRSlSLyfPedaRrAHZXI7vSeWu3EfRLjcN+3dAW
ymhsMjR0tbVBJe1/14+CFsTODtbPGpmcguDy+jAUTlBQmBjk4AZMllHfhPMpEifNpEwz+jsUkDh5
6vrWgYLcvgorfiq+nFvI+HOGLCM1aTCljAmFcFkGJ11SfAvhCcNOtm7NKyvUiwJeqeNQjcORKXqW
7gsnqAlSf889q8/rWtcn2s+XfkRxgiDE9lOuXFesf54980SJDtLj0txzNeqDXN3PiAFR4KjVz2UD
dnU5pvXeyOL9k2AbYSaJIHKyyaK/drMZiDTSWkKpATnknQotM69CwQTsAMhBAjbE0lAAnDrL8SPy
hulGZHv3Qp1/Yth//mSFICr/epOJuQQY1tdN1u0CdtyCUwjKP2FhnQF8Fuy7rX9YVz5EBMGGHSoL
CdGuxRB0UlovlUAXVQEK1sp3x08NC9QLM1uWqD30KUCng4WpLQk/1gRXIHi5IZsExwtQxvOFUdMh
LuFUxKLLT2ULJZtoXSow1n41Rg9Gan5kAJ4qbanwGXRbOPpyW4l4rxAfq7VhNudBaoRt7VAiEKqX
Gir6mz6LHUyQFpEsjLw2MDoz4BBkWPwdUvH6hzwU7iFmMy85udFIdkZXAKvfQxXw3RPLfxt6A0Ba
vWA3gt/4gbM8VqJ0+fyIF6NtfaBi+ClrcgsWsBT+/afdD/bwDzUSjXHup5UWKFIuUaWouHkZuSqs
snmVlXYGxMdqadsMkU0nc9TFO7LMkje5L1QNtK74T9w4FXRwTWb/L4uKKbgVU7NAYvZdqeKt15He
LRDxtVEfGUYYtvkxNr5t4MxjygXXVxnSCIFk8Hqwpe3fRw5Jl1xdE+QGGOKmHOgjPewFH7HYmG0J
E7ffxgZD4mnjx4PEJnGT5ZHArk4El1lvvUGJBgX1SZo13iD7K2iausCFOT3snGOhTZGuwy/zYyo4
WlqyY8xf2yMvje9Q7QMimONA63qIHOggLDa8k6QEAgvbbBKI5ui05myjGSnBS1v8jECQeSZ0MYqN
nrjGTIiy+U2i3Tge5k2ftMllV0uuZ+zHJBobEGOgMm+q7sSs0QL6GD/yfI88ISdyebGt9eWN4atx
B3fI5JIkYF4MZzEF/Mm2vqr+BgHHyBduhXy/XoTdmSzFj9f7NwoGBWhebwB6ieLL4pWjfLh2qSaQ
LwDeIihgtANG9ytV7nRt+2XCGiYb39wSifksOPGT/GPUNZVHLgp82LrUT8hI0oDQsk/zP4p2emsY
xM9jya54SinynJFIjl/MpMa4QoVtVNG8SwKGmBFyfEDTphlY0ysrplC0NBxXajTndWi8mD0Iqycz
QHzVgPsg+bWXkEED4iAbLUBFEM6kolBI1YFkgT1a6H0HL1TpLuExie29sEPyIZQ5tQ9O4bH3qYEh
hkluXPvxfQ5UybE+eKVH3GJU7IJg7W1Ga5ZD6WocZNr6HsRfRNxVAWnJIY1zvS7wRZEAe+b7x0Jz
yC/r5LzigaWRuK5vidbOvXizZZnzTbxONtq31aQ0Za4tZuObxpt9UldwMVvj6AY9o20CuXr50ksc
b9GhF1BHV0L9UaB89Mcfa+PTFm73xlyGOe6XbM3rbg3DuE9bwGprrFw6VVfyXa3paWuJPNVjXQLM
4SBNhsMOKbUMB2iN8Sd+MvXvSasPY0FgbqNtSr2EHDVSLRVJE5vVtJCJxz+WN3rpqq+2oFcGnNGX
LxmxiG8AH4aHQlq2/Sz7gds9MGRMrWOOOZpDIyh3upH+CTpsg73n84dlJGPqckwY8jIJxHtE3aY+
jFRWH9Mz4CHg8zyPtQgS1bN58NwH7VvoHpTOgV1SYa1oTTjH7MECV4ChgcBzp8D9Zcg14vttT84E
XlRAPMETo2xYKpJGX6eoPjXM48hZDj2G/zf3WDA9l74XvRimXZBXwyfCKEc1OByjNcGYlu+xHYx/
MmviumGL5YHIJYrtEGYF+XecEtUXrLyC2z5KNdCWN2dnPefAKebOQ6aVJou70N+5lMYNUnqjymEc
cWN7fj5uUGjrEZ2gE0/j2IG2oNqquw07cZw9CmsDmbcyRXp3QJNsK/ESN4fjMmLJ5vtGCCxCtTed
RVui1O1tRICj1cVvrHzGdk/BaTY6aRrWnE+HG3RmRMNFWs4tvGEhOQasztrR8kbtrei0Z5F2vwoF
tHgeyOWDeGXmTl4VrwvwzCr65RB985CD0QAhDSXarvK0Tl0p6eI1bvCa5HbaN7zSpZWrdA6rW1Z6
BCCGJ/0imp+LXFkBDKhGtEp3H1I66RMQp6b+UGX7dxpG5/onyVlHS+nCjnBUxQWTBQ2Cb1/TLRHe
7GKB0hEFjSg0BT73rdS4UcR1VXtN6QJNk3xzJJosZQ0Ia0OAPFa+/Nso3uVTfpMFljr7NlbpJd7K
RTuqA4DEWeqIbQGbBgeFr/y6JWhfoTHxc0kfsLGZcFjZ2dHhmN4xZUSAINczCL+KzG26DVTKGIH9
yqI1qW00z0ApjSlPVFZoN4mxMxrUsFZ5tnoH7lD2NGRq+5M9vUmYfm5P2tj0+Tg/NF34ErAf4am8
0r1eXQMU1uV3+J5rI2RBcwT+jsja0sWiq8ApwHEbzlEOIDiOTDRCoEJ5zqPr9x1uZTCljkFX9odZ
OXBWiIMXFTxF4xpUGa0UYSuYL4yGAamvwlh6iMZgkl9caI29f5GeO1sq7McTVNxiz8gm9JkTvSfz
cu2Zc0ck+a2xYzd4Dk45MtNUynAjJinHDhiRK4KlHbHwCWpYBSc7pY1/Xw1QdzaYXri1+yMNsatK
NTRMUD6vOIUFz5WinLayfio1wOszHCPjklixo57hoWaxCr6a+DRyi7Rb4Wg9l02F4i/+pHdr1u1F
VxvAEBDGpIzSW7WmuYU9S1aTsY2IbAxMwYyYpZZ/Ccj+LUYhhQeDoSfQpDcrJe8PNwHOkFN7ixoa
oQuCtrdd29wQogrq/I7NSR24ITX/ew+mxfB0eYW0bRDFYoKMA39jPSAeLjaIBeXUSiDbOudzVaNA
TjQXZJOcw6Qf6J5chqTlzzANxLsAWHbd9YSn0lqkcZLPqfx+wEWx5IDcDMX0hH2q/rq9eETQS3j6
IxU8yf2OcfLBNkwpavR3jexfrJnl1dlcZuhTxXIkFlR8Qx77PADnGX9hVstVObA+/PC8Ccy15NXG
cFtgt8f6Do7elnEG+ooDoUgxP/mQftbE6N5cr2iL8yMV253MqcLUezpXm5sBGvjRQnsmzYpqdFye
nXxSJ/sPzIl4D98BQwTX9dYgLlb8wB9rXE9NBqVsT5OQZi++KF3e/1RJS1kbDBGOoezt5bpPNxbE
JRMwUjfIAtcuEtkcqwzaH178kn7ToRJxwRs4nWIEszb6jvKoCU9Z8kLhY/XarimlsMrEZjjvza9e
DqOxmkSDwrvbm+DH3CSumAHvo4KskHXahI4NSfadjuOEX2DcTC/qcMqgL1dEXivX1u7R4mXS+YeZ
CdV/BnvMkrrZ0xZC6+oSHXhN7O3vWkZoDPz1dWnV6AIKSExvxHkT09ET149/O8V2w1eGY5EplFKH
4RwhLv89nw1wGb+n4nRrg8p2U4HwLJhiF8umk6B71k1TzlGSdOvzBNhPhtlVEcsun6HS9ZVRuNcB
Y0oL1akkaN3KPffkybQPi2PyIyF+v3zaBaEoBH5KbyCaKRWTlnEvVRQXr86eYfmC2hl7RWtz/ygF
3fVu0wvyNewe6clgxUc4KTUvtlKGVrXaHVWkts0ox/M09P20kAPDfZ3q7EUlrbAF505RQdJi6txh
1q1EAtf+5riykzHOzjU3V7UeyAQGJ82oAuR0+sbe1VOrzykZ5RPn7R5TRHeZQDDHN1MPfgV2+Plk
NhnwKklV4iA9Be61jDoe4iPA++xRU1U4UFyyw/SE9BixRIjQZ5Th2SwvSe5PTj0XoWRmpFFHR5FB
kn2I8AGow2ZEfdU/iatqf9yvzwZu8i9PVBkLg7PGlFq/1lj4mSNiCwODNE2xoBjtczrby0T3yj9E
+Fc7tyWYZP9rbVZOysvoeNjjCAfizB9Nv5Bma8laVlTkAQuymvl12tiAas2zuZ+wzODQvzMQDW4R
AN783x8oYQW+TgIVYdda0Oi6qF3hZaNBxpEieL0pV3wd5IMdWSXaFKXom/eFvd1imX59LVE91nJy
6ET7uRg66QAb8v/gyooTmy58X/UCgFsZNwbLA/MXA+EXJKSYpR/b0jmJdOP5wJXBhyCvnI0vXepA
7KAoWJaDRPcH5idVI3LIE9ddCntKPxUCpw2JnPoetwnmYHDwN/6t7+FTCvAeqoligpJdDzqhFYul
7C1QpWVevTWcputK+T+sgLvnfUfx8MBqKskQOfKKem0GH2lmGyYG0nXq4yg5oFFP54xdG7rEWkfI
urGYngTaoWTcmaIiJFCLIVB4vHXba721g+OLNOj5R0WdQeIfLpOfFVcrQ5lYYd/lN22MQMLsEBAv
DfWbl9scJ0HUphDMsajSo6cx6DG3nhwGep9l8Ehw24I8nO9lv3vHaPvbPM7nM5XdI3qBkByycm8V
HANHqy+jODNxZkOHWSB63ZDIni5ldgnktqd8/jzO7frkbcGcU+cvsAK9k6FD4eNQP9QhyeY4zXSB
VluMzitkgUw3xs3kXWgRF9VhL+/2gB2Imkj7BH8UfBqqKwFmTXxvF+DAWP7XS/DinZDGnqqGWyNr
Wwz1mdp0QX5mG8x5CTtqbaZ7McyyBSbwG/O1z5gNnNrLXIN/GPygXCDURoDhfVXZvv+rX2jT/9hj
A4MFGquoRY6pikpJ3wXcvMLRvnKKyVWX7Thz5TQsseyQ6fym/pndQ4Kg2/u7g81YURAHcz8ThNSC
9Mje/kWJRh64/f5iUbk+Nedn9QDmiH7mdXq1bbaQ1RPsfF/fGD0J9e7cGcnj9QXVeudSZhUToBNC
ahYslaaYAFTHWz+XY1gJORcy93VBtO8x3OJ68DfLV8oSXdnPt1xr2HYEfIQlGocNWJA2D/GtH7Sf
0DVJZUWTwsMCVlJBKVJEzqfkTQ6c67nwbFkzlbmn8Vhegs9u/Yj7RXFD2NHlbraORI3rmh5QlPOW
7g9umzPeKyB+fdsuqGB8DQdBKwLCrGzxjI4OMwYNpgP5vp0y+wqhwBvrY2z8wfbf7Zkwn3PfBQsf
4Iweya1bLYSNWZRwhZ63PaFJSkBn+JQ5rdKhCLNiYaLjs0yVLH6CajOYJzen/UA5M1wLiVjl+9Kp
oSbDdW470JnK+8Wniu+IdlbmCYf3U+OONEg8sLIfm7gBrwEZMS5LpVenhK9CSsTLSnepkifAyA5Q
1rwdO4C2vLdv7nLXwsdAhSN2b9+SWpjtwMp9EjENuhJ4H/7e56+ziCkLEjavgJQz9Uuj+NkAjL7O
2ICnTUdv259+2yXJc8A+Stdblj0Cd5v5tXgbgKMsBubMAIRONhQeiBpi1stvEPUpcnM+4A3Sw014
Sm1gmviQeV8+vX1VJGX5EYlikeBPpdUqfHHcUoyCHSkOtmwSgXLf+9KsdMC3LDKFnGwTqgeBth/U
5+pxHdkbjDrdzubqRAkeoIZT5yehGc58fCwbXYXlnabc+383T5KtkFTZrWWoFRal/iyD6hm1Hs8e
vRB52AkNdLaxkBO10AAqJQi2TSeKbv1DfauU8PRewiMa/AWOM9GY7qnNhxyUtGPDldBuSif7yRn3
YdXXtgg8FAcQQEe+GYXcQ8aiWxuPmbzTTevft9Z3MrEbpWJie2o66H8RFrhBW90srksSyBhneXUd
lCqrwhLiZl8liqAReWauwlFThMzdYR4kbOykCm3Q6gRS0FL9ggX4C8ijcjjY+ru/SFnf8eVngzPF
jlMPMoyBuF4LJje5Yg0uBm6L5t2Tp+W+khuYfqiHyKENzcjuCTGhzGQQ9TKtILFSZUHiVrCOPpNx
+FayIz2JEpfBJKqT2vWTN1FRBf+UM0ocvL2o8zaDZ4sai6Pr9I7c+pdteOouETgVuLobyeKoBSrD
x8BLfwEvgzc7xPiXZgSN/aUfI9rH9XbLR8WxgeqcNO53kYFVyl1n+AgYZysl6yNvwDQ3iaToak+8
UkPz8DBG4ksTWr1p3kg1sgtynMdxYEw7foY8m4Mz08L/p2DBhMciaNLAi/ZSA2yStcn73Y6DOe8K
p+UEPMbnziBK3K1Vp+3qSPu4MW+p/romKHmOMO2wb47n9drPcs8Kcm919hxcMqmENSPe55LaHTFu
MgSnw5nvatfdfjayZJnzq8jCueuDqMuFSFDMz+BcUOdydnuyJXKJ8oJQj0mlmF/ii7mo7QpSHGyp
msYIzIb49zU8qpS34tnVcUwTzLNoz6wVV92qazwFkRznL19XE3krUdDL7XLXq6uDRDRfo5OI7VFZ
Ky84f8zrV1tR3Z6HYAU8gxQj+/VXU9U7Seu7xiZiWqb0mf0pg4mX6p+SBrRPhV0kheUsaMSmVkJC
qM2zVcCLao4+Dv/ayYXRJrVzKxMfTnW4rW7J5JOYTGqQPPnwQXjdM04KTIWx2ILSBaAXYoDwl9TW
riGt8hIpsqr0Y5bADugPPZJZr2bPOjX6rmMdwBIrE5hbNYib7Wwl1Mu+8SciRBvY7Opek977w0JT
y8N4VQ02t8phSiplJEwNgPey5bCTbHDzCrKyM4ZBLus/igE9teXmQynOMk0/lYPmptrB+N2JsleA
HKef8eKASb8DC1fvJrjuwzeO8Wcdh4J5W7UG9OPZM2guiF7HBO4iT3EVhgj+ignU7z7oOgdHq9O9
x7cYzRAv1C8X50zWc1nWSjpWeSd6IU0EB/PK+nFkmfzTppxfZXJ7i5ZVLWBVV7TGNcg42HyPVyxh
GaRzNrSlgWRgu3v79oa5/f6zWNEzLtNpk6bblA1qNrUZ7Wu+yBcBqtv8wlpwoaZlsjoLKoNaDOSd
ZeHUFyC28NsqriW2gBhwwunCRivvn/7sjh8laMZCJWqVNOdT7c6RN3l7OeJf3gqsPIEhehIKfe6b
XgrtzsXl3SnNHPUO0q6JcC+X7iigE4OEWGjpV32fDGONvC/1vc7NiO151dx+oBdxpCLZJ9B4lkDh
9Tw9BtRVHLrrtUzQsTq2iraV3J8r4Ig3vYuhSfRY3qOj2M56rVLhBEnFCkzXzmJ0ur1uneS306ET
ONwSWloQRvzPrStRkpVCoVww4tjIsd+12xYBlYuF50UcJxi05K+zfl5V8csQNhCzskslq36KhP97
Ct8uwJICfR3Udaa9UgFC5lJodRpjj/8HyIuP8fd+U+UxLIZollAvcaeCjdsUU65qW48XZ+wKe1fI
cVabK9J2U+u0Pe2J/GS3YHRzZYXxw+PtD07BxefqE5rpvZOUHq9Mk2Xr17JnrXqlx0HHK4UbzQEu
JoUEqbJ49C+6OTXMwCCXq7fNwTkSC1+rjRzUenYLhYtNvxl1HRk4qd+zmQw477B2eT8JdgsodRVs
DZ9mAS6Kqtc3hOXO4jJ+bkZs4HCfhLZC8QVH8KfEnfngHX+7sy3aOZUQgyEw1sC5bec9ArmdOESU
XX28BgM26p7qmosUFN4ReU6We5lC21tKipcegJxfg5dj3yGs0wfyZhamQyFBuA/5TtnT00l00fGo
lvG036FEQaLliTdbLqzJ2kRVGDsAQ7ref8EFP2xudwkvjlHwKMsfYFhNLdonCpMLeF//L6ANWJHN
HWz2pdag0iPrb3Bbue8Ms6E03TA6DfLHr3nSsH4X5nnCyotj1/Rs0VSUITIsiZG2znbBnomixhrA
IdTwbV/k809fF0qCbooVHKCEeYpWdPmqa4cZ2tKyUbtnTnPzIrYdkAOtAM/kZYS1Dm6FzLcoCj6r
thfBiNPRW+4V+Z/DDqlKsb5N0cWHmrokpyaLLBYeGHqZj8Fai/FRd+l914GU1ztw4+VIO8vfXLcd
4Ps0XOi6Ju24ffPpgUhrNcAlTmUeA+0cukMgjHR2o1P1g/Yb7XzsyKs5uo8CbB77q+BHzlZGAlrA
XhZqNq0i2B2yWVU41aK0BOXgNzxE3g1HlQRHudIsVfN45hGQHS+rM6eIbi0QowLflEZ8QsYpWHnO
Qe6oUYnTi4P4/GW0SrRK3tgQplz1S8vhhyLgPa4ulaHWYaoTWr2KCDyc+sr5gBFdDDEROcIrpWdM
xTjGiT7kNTGupz8YIA36eOJFiPx5/ExhRjRJWc84CuHcqoTrEg0aybeesPhcQ+j2wKrRmMSzi9sx
bburlC4bUSkx6dJtLP4+qKLchEfYcjwZavbYkFXP2tSGdUlcA6c0hmmU5gomkH7G6gquWeTw751l
4oYs0m1xD74qiMbdo1aN4fVTIDBAjlTD9yFVHkcc33Bv8wAaoggAQ98M+hzEzS4GbGalTyPpXgL8
ke5pw+J61q3DMu8Da6FsP7T/uiMA5jKLznicpENP/37pULzzKf2AuwyARyJ1z7BCoNk+B1DdPIIv
9ElPRhEVgh9MwSTqS9TZTG75OrCSTRh5vEUzYq8W+aNM3QI5gVmCbi97McLq0hLsAsEnxlK8juO2
+C5qpopZnkLVM4YBwdn2885HMRZz4U5u7apAQfI0l3ubotPR6s0IH/pHW+yCKv3+ozn7KruRh9uc
FyIftjw6lRGtokBS7qjhB38LwHc8Y1FPWs5FoQWliD8KQUl21qWTA0LTYRwNPKTSKotGlPmTMfUo
GKOnR6o2Z9/ld3YDsGDtIh4MJHvmYlY5tF7RP0TjZ5uQ++rN3f6S+oDNWE3w31AtNOfitMgMWUXV
ij0y08Ay24AEEtq3gAll8tWRPw9+aqCvZT6F2fgda6ZSvO7XmEvaVj20WZn6Va7xGLYnSivOOiwD
kgwKnRALBg0N4wGkDlXRNFNmxDF5S9qNO3y0PHm1j5S8L87KKzLlXJsljWx3TE7pZKybySTBQTJi
Qz7mVCGGzBcpwtbCkb7n+uvpYWl22tXny3+vJbCRyXJFiGOGo2l/Vki2lMHMP1XXe5n1ZRoxgJmf
uTQWWS54b91vTBZg6V2Vgw5BksMRazqgINgkBT8mOEgbIo7macNQsjVOR4qtaxz4AuM/oiCowzSz
OtN2FWN5bYStg5CTPAacnCoNSd6x8eCB45Ynq8C/Hkq55cGok6NNNtyvIj/YBRG5pmD1ZglosL24
+BN1BK8gcsu9LUxdtknrKMwUnxTL2OiM09DkD+qYm/uF1TSeQseUPK9g3lxJORzBbvbYNzXY+IjH
LucxPCVY8h9BMLohMqwEENvqHx6jPQ/ire3SFAG1hC3sAGYD/XeJSRepcPskjHCoA7pn2W/CevRe
QsWlSEyg6bTnIIt07RDHMz4JZMKpxj//GhLKxje1SZAqSqjYaRMzxlyAKIgp0mRRySu3zTzQ/mbV
nWnPO6kJAzncp2mq8PZ+DLOuLtlGwAXtpeIeqflpVihT8wVgTQJ4xPFQfmBjk4gqHLHvLPBKKxdV
uxkJVv1JUQTeuiI9Tm3hXfm2RX+X5CD7G+pMw0Blsn4MjZWjEpvAOaXj8zehZuor0r/NnDK6ZOnm
4CYDqKEedvWfu5jLxpHYWUIcd+kH0rLZfqu3KMkZpJTQ/FOlKmA2AzlpqDe8PKZA/oga6v0b/Vst
7/AcmH5mWQkiPHc3TCJhHUlPac3F5JgUpQk7VtTTFPoUWgVqY/28NoMZAQIwzyzwk64Fv+NrkshY
hI2z9rXNmTzZBn8IVlG/ygfOMbl6pWEAhX3r5+zaXcqiUR1ZtiuQPpsUvw90FiPq4kgfWhR5lA6d
hOR08YjJTS9TVaQzLzgDXzxFroee+RlR887G6yFR+UQHbla1i8xwDQuc0NzU8Dxp0gVBb3uFhWf/
d1SpafMkyPtzY9aQJpjNz0BOKlbRoD0tDY3NN48mYTQcsAjfBg4tYw8heG9CBQcFkp5vOGWhy/Kp
H4a358A18GoXSevY74xpc+zMneS55RzjiHLVIhuGbmRQ4P6TezRfKw9bm9w8gM8NWiQoRAF6hI7x
oF4w1wwM7rl7RVmy294rF6yW0F6z4bpULbc/mWqRBVZ2B/Nsh+3MRgLb6U5q9iUtPL/ooDOhZDlr
bfOSk2sqRSfDuLV3RKqzikdZrWxYihAqbOORglCQYe88p/0y4Wfn9/ngC6VGzG4tyeoSQqIdZhdo
8EOhitQ/A3pg6f1h/fgnOTFKIcuVNwLBOJF+hAlVXiEo1Vv9SNwDjE7JxwtXyriiqbQJvOFsYgG+
WFf801KEPLQa9ZcjJav0lQB+S8o2IqlcCkwQgZoVvOTzXMie9IAg/RL386416y5jU4+vvNkrpxT0
egbEKvYORORvav7m1dAIxUZj0QZBKjhwEKdjm/XLXxS3KOJmIz1NRfY4T56hGFYLl/NtQWVuLS4t
RRoN+Sa2qtx3Y9/F5XBajDvQY/GA5fNSUytElSsGF35PxJVxd6jPGiwxAH/Br1dX9+DnNUm1MugO
6zCtnqP/8sC+Idb9LfVVSh5pH6P1o1p4tGvF84d+wvzq3LU+kJoRBMQvMVhzxxOUcBIRwvfLrNdj
LaiTehlKZTYw7EpMxELLO1CQijRhurDZTh96PxAgyi3V7TDP+WZSlhxqJA5TY+YvBfYNZTQHmX85
iTPzavbhrfItEoQTLEvxku9gzC2/+c0d8HwGPQ3MEa/FoGe1Sz7td3aTy93WbqkdX2r2oUgLJCPl
+mJSlP5RGYkAzOYNlwG96w87HM8DPu4HvdxMn1+hI6rgKW7RJ8DmVC7YsKRcDhODi9q4L688ocNW
IqM1ot4/EFYp3j2SwP4NBbV7hCoSpGk6MwUGAKtDg3/Ea5NcnlVAUwrvQhgM6xYXVORUOymyu7qw
L3BDEjfK/bgpBqwKXvBYcwfBKd2nAln+NOYMN3tTq4Tj4IlvvWouvG8z2lpdOa3v04VhE+XRESFT
uTkk3RlDmK73qgc5KEaABlSnRqBx3ie/g4uxNHwO/nejv2kf/JP8piUJaGYyOYwCWKv3wQ4PqHRf
6vxEFbCPZahr50S5Khi1VBLEwvT3DdxFDn003I10itntqgway5zgTI9qXLVFngSS8dQCCe9FNUWO
QOQNpDzMmv5qUjpVjM4yZurXVhvYI5kTzUsb7orhaxwPuyyvWmZfjcqV1/vJYRw5ZpW4H+QtwoR6
OIwOlYpXCio0NEtNSs5IRWGTheKrTdjbuKTdE5Q0Yj6YA4iFioTLSoqT/5cFHV8vjIHjAh2VbfZ9
XTPdpCyf72BolmjsM91dKwFPERglVYGWlLP9MfiuJcMqMMCdtEVDaAOH8jZJlY71Zb6GltJ5uaxy
Y/08FuJmluKXnuTvY5TdE102mb5Rbcxaub6KLs+/IuGb+7RxHJisVwKxdho/xQsBtDa4c3WaIWDZ
SfBjK4d6eE5Fu9I1vhT2XeBP0DyhLZ6+DgfmoVJlymTkUY0K0pS/+K/NSWeQpxVscb+yCSNXnrQ3
EFwLiqUVvMfmD9uZEgZggTEuEomAYrl+x0248fjiiW1zZE1Pj/RMYagzp/xN5i4TezJE9n1zZPuC
bT+1oHl+/pE6qYXkzG+uaI+qBkqDoAyHxcyZmz0lX7l1/0na7621kBa/ln3rspyIsYrQv7z6jgeB
8UDYFgDAwpvI44/yFp4/gPCjVrb6OvUPSVknjz6ueff3KPKQr9Tz2n9rudk984eTwDmM6k0tbdYS
qJZQgG7K0mFHfIrXKOIT9aX8GbrWiPdDaZ77QP8Ird8JqBCm34L+fC6buPsKch18DrIGEO/ZCHNO
JEnntvgdUs6BgXPy/+LIPC446PXqufbySgdFloW4T5CF6VslUv6klDt3Xv6BcArpB1E+aNaGY51n
Rwloq1ZqfY5HxqFa0LD/L0tHl3uRju6Zacd7k4x+/Zxr8RyyIGMcpXAJM0z2cKn1m0TIMKJn0KwZ
0iVzenLRLdjqoM3U2n1mDITIgBKGQKEo0sogdBgRn/9pNpY7VsIOINcrulVQWveqkVhSQJSEuGBV
HNl3IvAbSAcb1vxKaKhKiNwGC8rzQ7t38eskB5sl2aUCRGrPFrzRTibGA8e4vlRURp4hd3T3J9vg
SyrOMDkR/Lf/CTUrScWWfSarmqOk6Lx2L2P57cgMG5sbQrGW7hz9pZ/dWnlNTdInkO5nFUGTXh89
az7KPqoMA3SD7vpcwlv5n5DOGUbeLLute1ZsA7SsdxkrZ3oS9K8UqnKEmsWew5e3Q8xPtLqg2qgJ
VK3ag0QaDx8/4xHObG6SacN+yFg983SPw37EhGDyTGXu0c9PUichaMpBVnMvQ3xhYk/GkUXCDaeV
4ogTWgy9T1m1BzgoiC6JT+9vP6ORd969W7stzDZhOPNkJfoowOcEP4CQUKXDxiCRkqprXn4o5YxY
NsZyZF4oaHBDEDjcJGWx2/Fy/9eAsslaQNROZA2ud4nOy4OOC5GWpE5QLT/3wnU/PJ+uC+fKqSm7
kFXKUIYxN7k9k/mgI4Zlsf9d/kYHwo5CbJ0AzxdOkYlnEz0fCodxzq9NgmpGnRlFrKEsV5+y0Qw1
ZxZHmc1qUurPrn4deer48wZmEjFbagt20DxhxQJPAAOkzKp0Ydfyv7pDTLIiDtLTa3k+gK027IWW
om5+M2wj1ypjZjApO2nJ1LSGTftxK8+ryZPil2RrXkE6A5lmk/7Fo7uDLHOdFYpvqBNz3+VF2ZWa
ZDwiJhsRSk9J1IYPGTCIT/+biN9+wjUdd65AVPOVu2ht/YRRuXK1b5okjPbIEhG3iTijLdd2tHRf
JImLPkT7KYiZTUpYkDOJXrrUoZ3E9F1C/XOn0J5FPAEv7ifj4z+lb+pCC5ZHH+I9w77g5vzaP3iU
UkZXGEGINNHN8gHVZf7FaF9N1EOOx9P1tyggbxnC9M3yDRFtH0b0wALsLNcSmv2lblNo5Z1bipGE
g/B6p1jy1o1JMts8tosdK1+sguUnY/VuCJqHRfGxBZ5/UfMoTnWiEQqxafrI423Nh526DJcL+k4b
my/nd7FxKQRzJjgqc3ANrev7o//zp9kZ1hPUhRv41zphx9jelgvXjs++Xl/qvcLQolJCWQQmCoRn
tCLNqxIo2+gj81NcWzD3diyCewVxinbv2U9e0HHGBaGlePNzeXMkzvPbDVpGYg/SwQALV0xP94bY
W9j/FGJCTK2ipE0yE4JxoWVQ4IqjMZu/VJZkpZWhHa3oBjkpYmFozD9xzCWCYoVCzNR/8GHI2b4P
kLk1F8o/LgefOBcbFP9hGG/SrGPUZh1DWjjdxXeNg7Fw1RWL71JDZiDs4nBXbw63kdw/FZ0uO59B
t8djivEVOdQfFn9eVUlt2PnAjzKU4rYRrY+qWg4x/ZQX/6XXLZEs2i9nBVSp0/d3s9DhplxA5NV+
85M9yO0ItpUNwV+2ZCrr3WGrJf7nJotz0NtIXgBLm76g8g/0BP9NDq1Ck2+AhqGr0aWlf2R0WjtV
tRfLdegDBylAm2+qA1NS8BKyfXV25jkXuEyI4hf9UB5PtAuZYTyTfZqtQBjoUJDh9xLpLpOr5ZRo
4Is8vDN7eWPuynyZ30VYnBzr83+kHHsrW1DSt6RYnZP9F3G23IzQWscENh9UDc9S6GeTVVheDcIy
bciRb6M6ZDo9CTx59n974FBvmV9IsZdAmDFOWca4B+VsmFq50bJ2cc1VyxOXuNUJrm3W0r2kvopG
v5AhmuSfvQCRZbNjORMxOnnql1gy/759rTV7CWE4nFQVr6C2C6hqsNX2fRLN7Kr6ayKINOOVe3S4
PqmjTgvKSpC+7399Q+FdPOxH910WSRgr0Uea/IEIdZTW+QemKUSyy1mfDjUWzO7c5enTCgNAg8bl
ZC1XIch9xfxnUEBI324iVa18riZUlKYomFEJVL6COpgv5yiw1AnBOnWBVJL1RjrhmmzibOX64gOH
PxI749cKkLhWSfOB9Si1cGl/uNfmYNaLhxXCor6bx19OrT3KW1uKJSQ6jPmevgNWfndl44ogKvAL
kQUGlVxfwh/8Hr7oPUmLyyuGfMeqOTNAuLw/L0Yqiwi/FrB5PqUpiD2ihCG1DrL0sF8UYtggXGrH
ci0Sd/dfEUwBMHB0ucNp0Rl4mX98/9vkcnWFWStRwDhhr3WJ5hllPqcefd9RTSxkXEX4/xWc9OVO
Xk9jE843FuvedH7WXQuHZ+fmqx0F2a1SFAEIXzM4Gy3AfiwaS8utPTu5ZRIteeWqINdwMyL2FwYW
YmiTIZwXdAo0IqIj9S43yF54Lea7fpMjXJPyVRskfJij7F4ussZ4LuLDcMorva1ousMmKYqbZOVt
Lr72a+Ye9eeVA0MWTw92HcUkN2+uDhMLFPu7cbwjnaQ4/IDYnMsS/wYw+yEkxlRANs9QO/Nfa9ca
LgQxHnFXnIaE7XZ8hSVnoQn3ZBve+tiUpJwStmp9ftRhnUfHguvky1ThyJRsSCNnFjPbR6j0j7rE
qu/J5U5PSYy+VN/zW0Tl8Y6u7GorShl2wJK/zzXXUKM67/zg1JcOToIV0QGxRNUZMR0wGxSahWVQ
VYjXcktmI8IL1FThWv4dlY25DiLqIPL2n8NlA3SAjUGfPS/vXheihACXbmeE8jKuj/Guov8ulnqP
eEzIRqJx98ZGdZlud01Pp3ja9wlkNTJ844aPpckYuZfwTQV6U4qCtuH7gu+lVLEM4xc2/o5eR3V2
rLRVOuAInESNH6ypLuGyv4PMS0zL/MiuTsc6nGmc3C7U44r6GVEVSsK9xQTAG7K4nSNnngbcInDO
Vxy8qBX/dzVkz1zCZtW4/cR8M/EIRDvlTQksxKIoiazjexgMj0X4uNaa/VF/TlDvA+KAOX8mX2TP
YYBnIXXrog8a3ADnT4iEpvRmqP+1A0LCBvga21qukjBTiO0UVrqubXD/1vmfPPiwQBWPKk8dGJvr
J6Otrr86hN3QOeXbuFyoMx/2QFVUHDfpqyG1aONJpvMPyqpeL0PX1pGtjhLX634dV6EQzWILjnAh
3hqaGbGOTs9FRQaB+/W9qGor214NT710KvAkqb5t3HI0bbTnFwlExtWvNp8SGQvMF07UcJFiCQRH
EmER+w/GVsVR6nDuGRxLmIj56jKJrjKPQdac9uRyuHTZnGZwoAck3bTsDThQBsGuroqZbg9VkAKn
rs0mRjXpfpnrXtStjplv65+cv5KRpb/XKvLNpgAYKQPDS3jPKx2Oi0l8Nse+H7gkoyGa9z4EociI
maDwRsuWFOv0o1qBsV0NHBWJM8yqHiEWs6mLhIuIVVRJ3oOgS2AMIQKSH9dyNJnR4ptb07f+uXND
rzTvVaFM3ENWUjao61+g4iUAwfUwaq2RBSiLqHpwN490RXQmfJVIPWeRDZ6gtwDiEjp93ukjzXya
QZqK2pyi3T45LxKMlGPbLNOcBGjp0q5uhb0mXQCA/ppBsMqMlojma7Gs4hasWri1b0zLdfvzn9MF
lHzoV1vxK3oJgqcV4ni2o4PX1mViqrA0i3vZjaXUWXs0viWMXFP53mioGxAoIgOWxK/uDixaoLQZ
s0SHkG3Gg0KUP9Ept9/Q5vwsGoQ6bTbJ5OE53TiNSrgTH0i4oBwoFQCybPZfMaeUw/4arRopcw2o
lQ741dej3mEMhohme+yFzRzoq8Y+Lv+STlE31B/kJYE9GgrjFPaHknUPMwpJ0eTd9u5tY/Q+TZnu
ewkNQ3UiSAf09KaXvqm4nRT+iSsVDZlGzJ5HLa00NswrPMnBBtx/Ni22Xp1toR/XyuebglD2GwR+
/MF2O8Es9ie4mNcaaEjSsDHz7QKLBJ8sg1UvEk6mv7zoXGHCKBmQQCc0LwTHr34GiYEVdrjy/in1
IgUiemtJhWI+OvmbYbxjId5BgazDMY54ZrHooGe7yFeKkUEpM73B5EGJb/cLeOR51eaQJNiqGvfQ
0HNsqA3FhhJ2lLxl5+MYDUnWO9Lsc8TNILbfNiFokpLpZeCCQQx8fSy4oKI5P7Ia2rBTbENLHZpr
+Aj3I3yRiGeXYMCLKnuTbcCU1OV+ySlVwCY5ziYHuvDtQpjAjHHD6X1ATgrWvqi0YVJBwcK01gzp
zCO/+uHPisMg66uFsf4CnuRg3eTcNgDvQ7OBiQWRI2pWbYLCmN/7n8fXGTUJdNL/wpg/aiSNUYF2
udm/cetdd8EN74iheW3l2Criig8TxdeO+0Y6GrOh3Ak9w/Tk5TTeNDp2GEpAdqtr9rmrZEmeaYUA
9uQyTRxiQ/3i3s071eG3C/WWPtePThrdUuMruQFju0uwPxVV3mzVeYckjWHrlr87JeqUDPxLLHID
WgF7ipEvqjXMeyMIzhT+SdFtxp+rBqO8ssq/pa+lkKfIAenZYz4Z5PpvZnjyKhJj9gnyOUlAlCLu
V8ItA97owclS2BQeqLKGqgw/4i6+01ttbgfWuWwUcGfmkG/uGbtxifziSuSOlr/Ag8NKH7XgVJrg
ZLw64uUtWyRxykp83cAbcK704RdUf2nX5Bf6S9RCV5DR9V/AMl98AEOlHM3qKd9bneZoRQ8d0w83
pNZXBCTAppdK0bQ7lkojJyE3gaoyl2CUvyA1YIHxN6DOzVWAU+51+2rktb/LLGPugSGciG5XeFI6
OaBIsK6/llfAsFgLdUa/oxzgbkC5bdOfQQyECr2oLMAu5v4YO8WulSfJiFYnLm+d7WQ5Hs6CpwiH
RYSOBAKWkLr4LPHUo2TtQ2CsqKqMZ1SML+hD3hRk+TizrdQKRM/VGKOU+q/RWj2Q3XvVY6Jx2qHY
A4hMyH4xcmhcskHoEgDqlO1wCX0Ae0r5eUoRS1y2mxz+mntPuHvTer6fCoSksBHEQP/j9G23X33N
8EQB18PDXONRPGFvW9p2lmi9idHvisxoI79H8BvR9i+6b02xrjVbxc7x9j5tIdfkPC18/jEYnTyY
1LDC4s1bwPSXA+BNKtzU1/vMFmv2G5XlLxd3HCrEWAFnIXYfcLI78lri7ZGpZjlvGEZIR28iyjzx
twh/9qhuwFvv+X0uXpfMfrMLgsKHaJYo79QK94YD9fjnRkjWhhIcEStQC9h8MqP7d2g74LGZoZtO
R1BgTM6ZpJ9b5uCo4VIlTo35Ds78c1VmTR4PrEYe8glTQG86bcwKn2JoCWmELGv6g7QEqVcDPyi2
5lStXtRXFAqHnC3Tq5M/WXk6kN258Yrnw343zv9mpsaF/a/Zepd+5oMgZ+sjthLvoyMvpvyKaqTV
n6pU6aaY0C+zPiwnAmYxNjvQYEf1NO1JD0aHeqZafDZMwcHLeEaR3i3dlbuP2MGtVe2TL3awia2+
3aQHrtCDHLHTagnlvv95LLGL3icMTdFev4g6GDNTWpi0gEIB45iJcj2saEf6jilYBausDS+T7Gb4
tbLOTDsfinV3LnOsKeNQLuqnLIXdW0V8alGmC68PBbxv3JfN0Ok6C7KdgsBgMCStsyAIv5P4RHf2
ZKGrMbEtoqCnNqqro5/Q2jjTD+ZzJMqxw5icS8K4xJ7em7FUDguQJMLZlMlXCioJJK6JGz1wiwRS
UySRP7Opv5aUBlNYYaJC4upELWdORBMCrjlUJH4HVEDb79Ofz5lxpG4u/PEwx/e/F6mPpSYZXGpC
YfjwMppZ3L9EiVUFTYaac8oMXdvg91Epb56NAGzolk8Lk/bQKS8w56a0wFEzH2f21U6ejzpWvT/c
WUHKrGMPGY5cFi+g2yGzSVxzcFxVBwmjdrtv7jNYEX1HoDnYZIe4cy5hsz0TS5xi9+WKtNqtLWgD
OBxh9UfO4u/p9XQKntl32rM+jNcYZWbeSEp0vNmACFanUzGt/T+C/taz27Mo9sLhc4Q3fx7LCHn2
zvqYmnS+EgcRHChDtYp6EUFWJSJdkd+uuJzjcF3RXgK/lNUsR1bNbLjy/zsk4jRWQjY/rOV6j6/F
8UPrt27eG/3Sq7w3qmu7BFxi2EUlBoyrhjCdbsFb39WBFtD3dYkKXQDCTKJYM+tLkll1QCkAmSMm
rzlBRgEoI7Gr9ueQtDkWnT04A1AMgD7BzSU7fNzzwz7gM/lty9xTyrSoFR/XTk8AXt+4Rp8Oekxk
3s4YQC7FEA/xjJ7sIB74l9I54PSvO8U5rc3P36m6P4JQ8v3z0+7DDULGmzYf4YvTJACNXig4wM2y
g4WdsWu/xmS+anPetFt6ud86oFVf6R3ag7NKFWcc967dHGLfwOaDhrNzuA+OoC/STGKhyX8cUmKR
3RivC8TVYlVEZ4Tonh3afk3IiY6Yvj1NZ1NWfKD+jZaIFg56KOhJ/nHyqtlkyFds3azEq93EIfpo
D84x93sMyYYrxziSCoDaSXTahnkyunIMX0dug5SXcL+BlCttvTIjB+IyE+hs1hZ/7Gp1OZS1vxnP
EWOo2vgzcaJm3/jBd0rtN+SaSijSbOBGyp9bdLltFeVtSvuhrLi12uHIgrQZ6klNm3TmaudNILml
LZ4dzG8C5jAUDhb0ao2stq3UMbk1M6G6XlWlrKPaBnM24q/Rw1a+2hZ5C09ND6an+UNpe0Bjg44r
djb8jyW0faYJKsX/H34/yZcKRTvyeMT4MJc6fGf1FvPQss7qXKku0YeImGTiy4r5vNlwVQMt1p/O
A/aCDG6NX8G0xCO/geXC31ueWWbz21QkzvbAnb2AhciyhDgdODv/oj1reKMgh/uY/SXzv3w+HkNx
7zF72HcdHVUTvYztffZqi0h563fb/4bLQmLhLN4kdw6ajZsMu8nlglz8g4vzHb5OeJWQibQK++Pt
1G6I6PyXa10JNXbfXhZ5B+r9u+YyPRZYg21UULo8DxS0zHlRIg2dcdXlzE1VSchk+CuZmWAxNdJj
5wQEtyUEr88fxScAU1UK0YifonWI8vp5bqquXFebcuT6ncTo+YoitcnzcHiP7yZWXruZSpI+RUoH
zXHm088T+mYopsWXGrgnSQUzGT+vOL3Ihj3tuhL35RqHIEGibrPamv/v9eWise18DvB1oh82ro+f
307U7TlRO2HspVKPZeM8eoLiHrIfmFkA+ovHUme4selKq0DqZ2nHRa+oaeZY3CMeodHVEo3XDMml
UKcKjybEhqK4nngEUgCH0biWUSAx0Abby7boLVjNprwmg8YxMSEenLN8VtVgfffCAGvk1H54zHxO
OrDdaJQUjvNUftDj5lISigkIIVSXV+L2lf/XfiytAdtnZepXkrXCQKmvzFZky3XxHKwAzm6zkycl
ty5G+gl5KXgBotpEV8LQmu6IHNPDPX9b54VdrXnThynLO4qDztNfMeadJh4rb3YLgiBKRTVP9NFQ
MbtBFzfUjxu3Zj5liFejf0rFhg3Gl98KBbxidrRKTWXOE4bqD/rTehjCaN/zNvrdJjrqxZ/fba06
ltC5A/gTY65dI4UlUJfDIZdtHUqMWDzNtezOMZV6FH7tsw0dFfPvD2vMuSgyDUr7p35vkLeLrCim
pJ8IuHmqUFDhUMYNuhHXmyMtoie5Ri3/HGopSsGHyqr+iXJyWIl+yKGJKFUxOCqWQtx4du6rL8Le
X6CE7XI6puIk/3AB0+stHidf4TlP0cxei0lxPy2I1BA9WZBs8/wxriH0iZCj/eF/Xe1YPC7vvXSm
1ddPDwIVdbVSHRcrCnt4IBWfnseYXOXvXHFUjt59UDANo6PGUxsskdQaquyRHtiy+J6IA15cot1e
VZHbMipL+E21f+kLZX9m7IcUTusXaVHbecwBeMM5N0b3rbC8yuXGjMAPAg+G/g1NOhRUMx4ooriT
fWEIIT9likPBZK8BxXGNqPCRgeG3aW6IXQLwhw5HqiSb4DhZ7nj1ID0jCZUUY81S2kTqb0EaLkcc
yIOXmSfvvSWJH8Jwf0Qv/FjmlIw9FxzINkr8ybD6sOjkT9vBFV48BFOKwaMoyJRBB05SGGIVA727
sdXncqMU+RXddZxbw3WWIT2AZJhSja0KsDez7SQk7q+mcTjCMnkb3KVobCp4E2lDr2JPsUm+LzwS
L8YlEBLHotsd1/F8pbKZrzz1YJNmGDowX0idDIrjqq+d+TQxS/Oz9w+ijDx+QFAs60qlkNrPi+0n
v4B0rAQBJpAYeuJZvJ8nyl/WdHZFEq2QdiSRc+QQk/k8ysu00PIgfyegpsXjp0gTDytK/v5MIFPc
0C0mJca+I0tPJVC8PAdbrXHBfvlTn3uZZQfGEdPiN1Gdg/17TcOQZQ+ny6XSDTmjA87aBzm9natc
nd8jDgwx2ubWNG+in838DhuubHVEn+owu9swMDctbZ9ceMi6lGaKlWmxOh70ulKbZp7mUdKEMwTH
wOSAyC2iekDK+IGLhBYhNP+2MRZHtU25CkCEo3sBUuFe9Q40hO7qDFFLFb7zT+vUcIL7F7Uwnamj
P/45jjny03DikVK0+oHBdTBJkj20vDbcz5BzPon+A/vMjd2plMjNbRSik0IlFCkoKBAt6LKDIU+S
efNI2TqjJ6ssnJTeZr02p6RBCY1bOuEdqSbCHd0P/p+EGOHCKmHx85veCvWBk03/+bCU7JwPrY9m
vtEg+7tP1nocRA7zaD17TC9QlLyqFvPLArset9lsqk2C38OpNuKbyChlWldD9KC/A51YuE1youv6
jdSr69TAPI8p3Z5GoiOUAGNvf05KkMX/LV28hPTBI5MzHEvqQ2SkqMj6UeDw+EB9AfG9hRD0A3EP
eXwoK1fFI+hp3tQS5KAwYwOkj3v8R9Y4qifwJ3m6XztS2iwuwaIkSEc8XwYHwRFcm1g3yM+3XWLB
XGSwgrsbPFnv13tE1UrkSWeJfNP2KMk5yjpcrGgF4ZF1yrBfkaciuVLjK/ezcg3V9Oem/V3/8pHN
udeCyBvqUSBDOI4tI/cwN40ws3aWO8w77SztmGwdstjZZpSkmbFSVRw7G5zKnTDEVcFGlW8Z0XTr
pJg+oDoEFv3oYhBNwFeiSLP6AOw5GXh+GA5qk8cBPKT/kiOR2ZqCen+HlIQCyX+TaUs+CO7yW0Pz
KUGNa3TyoXnmcKTNbr3BZyiYwVYP+CXqv57RlHDjDPlOsH3EgJWqh/X1tOH3NwpOn+6PTVAGHF8X
4XYb1bxsS5a+PA2BIgW4OOWqFzTpcc4Zu5XhDK/NVficIMZC6ak7b6ytecvoK6BjjYOTOq/RAAF+
CX9KZdh2oBYRPxqgUBTeydkIXb+taoaJx07671lQ3Cieg+T4XZFZBFa5QwNx7g7FlNiRH4X0xaE8
Y7ZdQSabet1X54aiKqi3M6x5LAI67tasLkJAfk2QGrz6/NOA6UfhBHXKLazIYBcT/QzSO3+EX0Cb
r2+UwjSHTKwcsveeWu8ZEcvzmOjdzdw2+/TWqxceViHTsuPhxIdXg7dRHtUy+VAajkzLTl7ErLRf
/m5atMWbl+ixzkER51PmxyzeFEZ/k0bDtGIIxZlkeTKmZZ5U7OvsdTQxlCMJEhoKoW0BC/lsv9ya
EZFEQUctDcBfLV0d7X6jaXPyXeUKu2TC9VN9aw68Q25osx0j+x1M0ppkBA24KGO9Vgbgk+7t+2gY
IKfeDfT2JXhacrJiEnWRrEMIccQZR41js6Hlwzxjfy9lVwFftBKpAeKVNBAxWEmBIJFRmh0Y3ZfA
A2sOrntyItSEfakbRn0hZS/cWsRgqj5FKJiUUrF7jFBe28pOHXQbG4Xem8UgmYphPMf1w4b/Yf6V
UvKjhUVFO4eorGyzwrVvDJ7/SfZiqJhxR1tBhPN7h07jKjPTbfrxn6xivyyyDZt57L13pqwP/iaK
yRa4ZImCENN8MX6/5pR49umDgJoqX7th4/zd2ZXIJgg3vuUFd2VNplrRqKPu8YXMwzcPlC+06JuK
xtXT35kPHTJuJp5WIFxdqw4qRj+c8sMZgr60DzJoDdX32xB6tsRTeNucPIAY6Xz7Ic4R7lmddIuU
9efi41LtuTPI4od7rG6r6n3kOzqjuUcVsgm37E/PxLtfsRdZaJnlNnfxLgIrpYg7pCG/4yHbd0wn
b6YGss2AHCY5PohB4Gpb3JlU8wbFsTfzRVjVPjK0iFq9EXqBF5B6JLwmMEBTvWVOA9jpd+jYO/2o
ej0ciUMLlOgK6JRFpT4ILiQvAjwsxH7C2trMxgDZSkMzqTzmbeNfbGmyNbBCwDKs71p8k0wJArSW
ZEzoKgxG5bsNr1XqRE7ZP0vIr+4el2KUMB5nhrJzz2CbkQkMpibLh+GOJDSs6CrWqmroi0n1i8sv
9fQS/o7WCtj2U+CRjPtSwhsFZYglpaYotnw+44yChiby5PdtGsz6ORdW+i3fymvEovIUqq1X3VpY
9T71u+rslgRRk1Whe4xlRAyXK0WX1/NTVHLmZYVUGeJIv6OkwmQN7BOuIzLRDWU4xh2PwQoi9Rmi
jJbx6TcX75p3+AxzIHeMQCPn13JbPMcWQ3kyVcD5v/4oKIp6c7usdiVEKFniRZtC3ZlNcgN15fGp
RTXFaNG216LVSamgWJ3/AG9AOn+9s2yLBI9JuzdRDnEB2jvNkZwUsReQ3VKO5SOgiL8XVHNqNPny
0n6vbkHmEl8/e0UaIPTYKuWUnlOLGErhBbaV5CqdB5d9+dZBI7zFOaGjUGHoje2pLhpOvkldbGt1
d5hxyYrkKJXk+tZjTbgwd2yYdkbibo6WV/3m5lQ7hSfqFMqNYlSq42DIk3buLAs47WlbNFjAjWhM
7aJZafNv+9AAitqZ+q4cGnvzlT6kHhNzw2Y4M9bQ1oY1ZKGwpfP+TuBLmdr+cDWvqRJLeU3pIN9a
4dnl5+IecA1sFrp0vf+F5xOwn3GFYcxsP8l5A8D/b52K9KaPVVcgDAUrXyxMOOTzrro+m8ZdgyAA
ndKwM8HqZtAFRKaJQh++oXyPFcb0fLsDdrZ8orTPai62KvwjjCPyZJM+aIREcJ5Qj8kXNFDxCUGL
FsUWZjJ8Zj6FB/ghYHilCzsxQXGymoBXL/C4NVSJLH2wmRTzi/KJFa2tpCQOY8yohiNkuOBqG0cG
FZy4IaxLMhowab+62coe5CvUZSPYad+ZFHdQ90IQd4sOqtubC5ljahHxtUShVglBqEp2CJ1AYpy6
blpjmr9OMS5rY/xDkdi/E7c6bPOGPbl2D2w3xzi3PrVOw07RmfkXSu9XQdTyZkfqm0Z+wNKG/SBt
fqHjVdiNOqkm/QhU6m+z1nptSgihqvF0+S4BB5l0KB0n1qSpolcdOXKsD3jcEb7gQ1QETMGX1nFB
vnMD80Gl5RpE5gGnO31HVuBLywx+RiUXaR6XVdsAzmcp9eI8P9WSAf59D7Guc7HpKf58aTcYlYE5
/yBL6FxPt9+JZScGIri5sDWLGNgHWqOY8FI+I2y95vHttT2H1f9OVl5k4ApVAcXzI5hjDTkv4rpC
z5aORRmLR7lk3xOHTzE1juk3lKaNur0/srcSn0iFs/7H7pqDeOnh7INl7z1Etjd6lhW97dAftfIC
HcsBv0SvBZHUGXWmfzJtPNm5lm1JYYF/5DaJ+pWbxmpctiT0VRTTM34+ujQBDBKeDUWz0MR/Mj98
TZfMmGLKACCx2QyfMnohMxrb8YbvZQN7ldur1eB4QyLp2F4u4+BOn2VQ1wZmyJHsqFvLr6WGfhRG
xbRv/jfrTZ9M3tY5gwM2LoTDKfU20YynCXibL4r3il/PV1fVZTEkKybj5z2DwN6eMKCpfsVGOIul
gbIgMSdMuAjEXyhWL74GFo4eB08Ty5CRSZrOutQHxqLuwxivwRGDt3ptb9xi0kzrQ4rAqPNJDg/U
gHmD7rvVWuu2YIrSMglinsV9VS6/G9UCOkZ/6pzcmVv29vrkoAcl3/c6pyUasnJII3FCt3eItpYR
5SJJy9B/QQID/GShoK5zZLpfABGVGJRqPO6NR3+iYa1hC+pQk1TDWv2G2ZfrweFC6Z+RgaxBDbsK
Bg6WDiM6CbugTSrWEYnNcKkof0YT7usrK2JQGrawjHEcunYegpehSM+NvWZGJCbesdiJ2QtxUGeC
lPl3Olb5uzq8UFNebOnJULudjjWocjQSO/gAULpD4MQ8TM8cqf+QaBpHT8RkEAl0JiPgqiiL4ABf
/FOOGmVM51L2hJPrMDt06VLDUevhqUMA9QeQ85I04M1slwtp9OLFOsgxx+0aZ98665XgScPRl0NI
0XRdhjB8NhYj+NbPOVZVINlFe2899sSK4nbEJZy33yhL8yCy05P3UAI9b/Icx5lyBYgcVcd9AxdP
+JFeYS3hWLR3WRJKolSXRE6i+Fivaaaf0jvUudgIqo3VcwKwCydY7MXBHbEiEQdWtRejZ7aLSUw+
ZEXwCqVAvlW5Ckque+g2EK2n/i21abUmVZvuXLrVneCz0u7fsTx4f2v9kxvrp4n7S6oPoHzVmVZt
HeZSP/s8zEDUQXqjU1bDDhi/pDdLEbs4oiZOWlQCyQsEzwuU39rB2ylqhDZ+8jaATXiFkZICkYoo
VWyincKf2r3dv8AP60BaZSWdZHm/jWq1Z+BGltRaMfQj/5j72jJ6nei2WxsCV8nfKvqcMKTy4zIn
6VWax0xbJhVdDihVyLFr8VJ3Fv39CmD3tgnwqPZB/x/Tsww/yqYZYVvPYTgVKOnAbS3esvOdS5Qk
6QTMo+QvloTgFCIFyCgBhYqZo8n82zQjSkTpMxbaEySdlvjmc0tYxIwgghoqJKZ9ckvSffZZUx8t
H/x0o+k6QsW19VOCmoyqCWioZ7aB8D8u7L3tjZajd8MeLpjgiAwNKDBK70OjK/lQuks5QMuYXl/s
kYMx3WV2yJvONbU6q6XVyy5GR3KUzqWssEjGEvCCOwouOpgc6q4priC9quTHdjc6bCnPvYJdP5ur
HNJII1cJE4ow4E2dQxisikQYQRh+fFZR+QG9hB/fTw6sIFxFjYLUlBAjA+YUCpJr/uL2GDZ59wbP
/FMxTUXfNwLVMWCjuXoll1mtpzBBo1E4YddWUUMk+++41R0PBqT/NvPt6H3HORIUMQyGs1wIRj+J
/uFbjNrH9n/a7v7zVvr/GHJKrg+mzuEF544jrYjPOVVlGsZ3xxMk9a8WjHXrdbQJ3R5UW069Pqz7
g8PxN5Pn88+3XsB0aEbfmkFuvFDuCt4maHk5Smfa0a2Vw+GoiPzo8PbnlNpfhXcGsqG3HCNWFt+8
ztrZ/C5zU9B1hL7KPAQMzVDY/pxTaMWJyQDhFTYOm3pboqk01Vgjz0I/p1IxRJqjDZBbyrtXhVfJ
CBrUh4qj0OzHf5DF4wFykhj8/zklqadX9egQxrl4lLvnikYcvVnpSYLYTiKOuWPILIIqG/9stuWb
QabatP2SLN+Q7X9rYDHmtGMnNoKGchCE8NNUs44gRr51a5RL3kbrc1lLUVPr60pE6KusjM48m6iP
RZChuJOuzv8xRKnKvFq6EilXzVgFSlRIOvVn3rSidmlhroiog8vK2/ufJEZZOB2llsnG3lBeP7XY
ZHevBkdyQAk1ykszxw/Pr0UJank5l6lC4XCMJxv598Zx9rCNx9BBajdNHbe2Hax0Uya1XctN3xWR
HhxUhtmld4hOMaNA+sbKgDfe5JEaEizXVTVhevMXbnziONR6JRMe47bUM/29KhVUK8fZABC438d+
d7VMSvCLIhOicMWY7BXaCEbchye1aYdaBpjO4HCQdGeQJXEz6gDoKPOA+9jK0lH1Wh2qxclN8Uhj
m/g6RtmPCuRbHugWsUDh34Cswgr5rIwgSbqKPE+3ZwI/K/yYf+2G3WXrCxBlbM/chWfLN2vuvv0v
bnOA23vrFj6DOYWgXGlzVYoAxsaZXpRC/gADeNtkPoFycgJlEtALDLNRZj5XyhVNiKkZaaFDER4q
qPQxy3WYjqCulHOwU9PH9Gz/O7duwNSaBncbtvR448ELBQW+JSginDGsyXBRRZW5VH/TpOWpVioq
jGc+We6Ugs6a1KGHbXOViZ9g/WJCtQKH8wvZ+IExINr5pmcpNjiwgev7Mi8MIS98/egswDfbBWC0
eK0+CW0Qikp8VLKSXdHdc7JzPojW2BOmvBOthuwh50U/Zi6ZPYAdcOi4TaMAV+z/f8P1l39/ONSz
C1oRa0ywjPvBelP3TW1JMiePx1x22KsTw3byWrnyw5d1Fg2g/aBdgIqEmU+pzgfvqin/fJS9ujj4
/Mp9VbzljDtHgwoInMtoh0uTtu4TljO402AXasmVnL6ehqvzJzXuJovcZUCvRXFJVOVja84tSibP
+8z0PZAghNLaWhZdtIH3+HECljmdZvq28+Bn7kqOD1xeStcP4WZwgydZ3wgSlznDslLwD5w2oPrr
+UIrV7VoHCqPC3I72MBhSU+VrM9FSe0fBSCsVEFu+W+RSJOlCHGRkuvXLtDMxjDRjwM7hp/8hoLZ
B/WyYQBQUAy0Y1aM5DLH/Toaasmrcp7E6fcjtRWWsE7HTqRd5JbBsqRFXKB0SxP5LAW5Of6MsXyY
yov2d2miLiDhGUzktAXeS8Y75nQuuZFY6VUhFe7uy4xzeTNPRk0JcNW8c2AyhpBqXcOaohmX3/Om
bVb8qQBoJh1hitZsDdCPiuySJklys1UDRK5uFyaH4TXNGyUAZv8mWqHB/LaWjyf+j4Wf0/80+8x3
2sl2jqgLkBUsaqWVFPG0JJwEhoAqbDyM8ZsvOiZ5boXo6gn1QbRDJ1LhdveHodPOvm2vVk3Lifjl
R90CXWXX8ex+AtcrSIILojODI/rhCK8ZXJTH4ghHMntLrX9NUx01R3+fPuyrq1bIEtaqcs4wN4V+
L+OJ1pn70YMF7ogaV+fURycE0bDR2zLsJB9VBi4lt6b4pgQ+FmepsM1FAebhCLZile77GXVG0m7U
LTRlL2cOGhb9nDWvapdjjdlxZQDwqtP0kxjhO9OTAYqgVoHF/9ntLgQZkGOW7xx4/6H6KABd4/O2
7sMXslbFiWEofUeE52oTe7GoZv000Fhc6mOdFpp4AiZ9WY7/ZbROz3Hrun5DPSzqT7BtIAIzIJxe
2KKCK17TMlb/sMdomXBjuCRzjTfZOrA36ivNi6uD0OR3AkFK5c/QRsdrFRo1CZdO0i6e8YWyqNkg
klHaFgmCgY+OTFpKeaoctlMcnEqytN+FcIqm/bC423xvtE7fZ2/5kN+aHipnlwNP59V7YsmABqAp
Iyviz4X+5qB4TBqack+hIwgr3p3gPOkd/8Sir9XiSJm7PetdfWlEq0b8UL/+9TPRlG2kqjhL1T3P
QJUpltOfJpXp2Mo11ybx+s/N/SYkjStuamOClIl5u+zTkzuVNcc1wAgYzFyh96HYoQJhhVrkh0vN
FMwCmWzxiTC0uYqLGrWXQ3vUTsJd4aYplXlFus8fBFGoDu0+6MzojwFYq6nYDkDID2r0arRCu12b
atu0qBJCHFKHTHTurf/BlxpQgkHB70QLrsaWMfSRrjSAt/rfjEJZ/azq2BAZphgiSax76Vm8vle0
+8CLtfmX3ytG2p7+RqzK3gZhObmQek96c7eOQYTmN+chi45TuKh6xckiv9L3yOwaAL7XiR1pBsvA
uaaTu8/ri9uCtah/JNXibhP6PDEjC+xi8q4+67uzGWJ5wSdijpqK1FjRAQp1YOWIJSHYdnumOdP/
Y+3iPXSntsVAezzQ8000+nSi141rq/h/AtITftcdvXsiuDxIsiETPtqBTIEm4OgAcfGdpD1hQ8zv
17/UCBHL1H3I45iwdxWjumePz270Vqy+MICa/acpS2aEaxwlIMtlfqrOEUYzPQg4TNclSkygmv1/
z94aIMIf3rF9XhYZAn++pUp6AnjXxJaTYdRiYMQlZLpYLGEXQ5gqH4jmcUN/+LivycNKJ/PNK+YW
2Gfkp3rVKM0uQm834fS1XkCzJqXIBkHO0vVMmzLQtGabFU1DZ11i7+3ktr5m+BYpA+lNAWxN5aob
MHlgpkDCxju8H5HRbSoKClVWnpdxNWijsVD5A6fgaUe0n7+RYIrMnvmeIWhuFIcTslpokZ03jwxX
wrBDkGUq1idLL0C36M3oJHgTV3m46YY6SeX7f4i3XD7VGzveqNpIGXJJ5WiUoDkCkqh1suvqegCx
/kYb1mI7RgzDI8gxB6dyjSO/BkrDefSC+VlP7Ajy5ooNt0xssycWqkgnFc3ot2HODVB7i+yP68VO
dZAhOJCZywX+YhttlI1V5hgSqzi6A7+PjQ8TGPDn5Rf/CvFMxeMIFh76I572ASizuY3gEY+qau1H
UO4Ew8FuKfizPh/VfFfVZ/AS28QkABYnxnDn5cizDcKFo90peVw4l/OdscS4bEpMOYNFKVQPcnNA
nXodiDEaon+KadNUyRwkRqGP6Ax0e4yZkjSX/Zmd33Yb0u9iXjXxCTPZYGEVg61U6WYLluHKTSPm
mjCyCJYik8nvl7mD3lsKglAd5pd0R2q6M8QUwZEBrY3oDLqVjhuy962OTifD8U8hCqIJiizLLqwP
FMVbKWYb2qEeIRamroO/5/+MGGV//3ZXNK2Tq8zTr+CWYnHc+B3Vrx29clBhsjANY4tvzsRJd6ZZ
qhxDK18lQG00kxn1h3LfM4DqKr5q8pO74hUj2gNmtO4duS11lJI3UpZakAP76g3mxXXlWatYM5Rh
DWa7zWLcxCU9oFR02kp4H3MvH2USXyx5M2Y1eA1SEXCkt4AmqvAren678urUMA/WkCmw0cvTgeUv
2fY+dy66t6bkIPVrKaLYQUr0D8eU+A7ynHkuhxXacHo5zglyiZ2o9AqgxOAJL1HV9DtXICxQxtb4
nV59dOiP1OzcAv/R1OJfp10AWGRB1Bo/v9Hkic9TVUA3ZTMYzmfzVVX4kJLcxuBAgqjLJ/QD3GRj
9IxOS2FLOOCY9HzXFO0Tmc30GRposJbCSphTXYy7OuSeDav1hOKIahS0vcLNt6BVkYkOZvXBPjQ3
oJHXIJs+F77gUoYBGYA5d6lyFRjOtsUYVZ+G3HPPF4s4zl/oXGwrlWJNGRdCz2Vun3yZGy8J7nDG
+kF4Vng8f4dn0vTdy9Tglj/GMDu0KI6PrWtueu6oyOjvY9Pjt4nhozaxmOvBCGSx+9RegWDdz700
33722SeeUPCvFtr/h5ZB2ZH1o2MZICM4D2XCiEXUU28xE2AloknwMQIYqotmVEETP5TuyQVlpBu6
h1mhUPtsykNU7J5Mp/X9GHni08PFP4p/r2mtb3IWTUC11mmOh8c/BXCuk4Vd3e1jj/vegQgPlC5V
qrHQZwHEij69KwlHQU1y0ZZOOstcKQXWYrNZDfTlWG07KntI5VKW6BaWrqLqlrPFVi3M6gDmcWSV
TcepsRR5azf0b6kDnO2D1KEcL/laszFmpuHYVc0WGWMoMiud9hT10xJjDK1GARoJoSIG8Zqi6fou
QGgPaqeE5tDY94JnyKXNlI6alMgWTidt3B2WM4cJ2m/VCK2Xe9gE8kHUK/GWqlIbt9X7VCvrWg3J
wT6PVzD11Fydp/TCCCdEh3TFzPE9lxGvHatY1jTkLNTGViKZbuiPqRX8MbTtQ5rCxKCmknKg2WR0
Xbg01dEU3zFN/RDI3pIcs7lO3K9u+kLEVYmglG4/hcqpvFFog0ZqmWFMPg9J2pBKhC7eioQDLxUN
Dw2lIJzkq8ztS8RmN8jmeSMgD/fdXnJcBul+enL2fb21A4NOdSmdr2LzsoFtcHc12Qwpu/p83uqL
Lv/fpCqHI3kvaAg5jpQmD0E3f3jDdhx92CjgtkDsFR8ms6n3mAEZz5QNMjSiMyc7Zzjw7EALXsfq
8+LqM7RZS1At+nL3eeM9nUAhQAe/hqf33iroiVono/EYVC3Ul23lblLow74Adlxo+Dgh046n6k+I
ulXNklAmiaee1zWZnbZ0K8dBuFP+QAFDv7DJ1xOa5ZGsHzGNDuLwv3E2PUatE3e+mIxEQuJiaaK5
dv02IojaqSFIXje2pUqDtePCsKAZRABlZpkJ4Vbfjt4mCoLKimc1X6ASsX5suIP7bh3h/jHNnDSx
BNX9lbyfULjR1RJZItonbQYpdDwzOUvuzQZwup7r64CWYC1vjXH2SYIatdoWYuf7mUxcOD9keQca
WVsvZiIjw43BmzWIIGyUsvy91Z29aYSJy7tg1hdRBMcQux5lKWqxlTvnixZvEWeu+mCTG9Ncahnw
fa7Vy90qYWDYsVExY+ljfRv4zGM2YWcNdldi9Ggnahac1xo9FrCY2/NQhVv/64FSeur3Xcv2yGpJ
ob+KN7hGhWb6aaUkjhk+zlK6Kkzs1LpAotIvEidci1+tr71dtNGmhfiwPnRPttfwxQsAsKPCrm6A
cwRENzuf7khr/ljxabqXyvbMJ0+fsCX5k2XgY+PgSalBQslbeCByw/5fqv9yvkAAOsV3X8TboIRR
uZLcyR6JGrTEubYUx9HkTmRpsesVJ7/c4csT+tWpBcrZxaHbbeTBhqWU+dFSM2S6KNtUx+Ls/pk6
pts+Wm/sbsEkkbfZPbzdHzC4bhmq+0BTQLxG5MJU+jPYDGlaMY9ZYtnu3i/qb8PuS2IQuCoSC2+b
7L19trgtju+HUd40RgHFC6vUjhtidcRjDtNxUBLA2pV60OftRwtnFI/0woppe/uSE8o95dPT3QTp
rJUO0vtZp8J9UEzOMyjoOQnwPXk+1T4W0t+mvb4AgV8pUkHwq2JNkHf0Xu880TmwSoaiKdPPbwi1
xVyUvbQeqEBXvWCSEVlgxaIgewWhL141EXhTEKnm9m1oQTlQyIY6Y7u+WQX+uqhE2En72m2yoqFz
mYI3hA9uCvw9GmJACruthVTvtvJPtfrB9qrHmngu3nEg3CkOG2ax3lNv0q5YKK29KEtGRT9guset
58rSwf5Z8gSUbsfOQrXX3Y/JwhA1MXxqvNLIfABkq4maGrTpgv4a4H5mVRgWQ98QJ/xo/sqjni1F
6XJI1io11kvaN8clI8bWtWQeD6p2Jm0xHk6tM/8ngzCIt0Urljdwi+1z5JpA6upNtVk1J2MOb37k
4qb3miQ9U+Zrn0Wnt/lkUfqRUISAVKzNcxWzYUc4bL4I5ZO6UpLPG6PPQ8fHsoEZGLSEdayLKoYm
NwHG9gCO386BKHmYYzUyQLBkqCRAJYFlKXif8LviK7Gwyvp2TSxKe6QDAw5jzAIR9zEW4+ZyYY2S
DeUUkMqgqpqzVkwESlvdOw9Tg7HewXMosXk4ioVmjI1PsIUmPINaj0/Iac3JBgED1hBTPsnqY4SN
l1MBztX9pziDC95ItriBFMFW/4UKL7zAhyoDJWbHi7SuTdrGNEk7+FFbyALwO3u6fovpLRuKdraB
kZ5gfr3bLKYBPZo4gcBNqzRirHpiSfR/aGOv0s+PXM62XSMwQldBVKARFNYyQR1p9VZc3v0RioV2
1JmQ3F8J5ioIpYV/gTomG2ihrmO1IKm1+CpDdMz/RHMoVFKpXc8n12c5Eov+b4oaeudhdG3nubyJ
bF7Dl8RiYeLFG9xysqlRHLcPhKwa9dnTh8wED2+i3tMpvq46mVjaMrT2mGsvSfSlxfn+QmgvUr0Q
nadjqhzZbKedmNok/NrU5qH1xpMY3z+AqoaElcJ2cwVP+KH2Tz3gtu3i3aCJaH+QhA53shYOlXhh
bazvL0phRyLpszOJLodlEw4n186dDv3qL7rTjFqGZ3Qmzg0C67S2bUHElKAmQd+6U/FroRhu8xmR
2YoFmC/sSNaKnivU4D7M5O78ev7tkyiG/K1+k2HixSzP6zKwWOIKXhmFQtQDrFcv5otO4NggO7Y8
YO9lkEzMZl43JQ1RboU82+KldKtVdan1lTB867obSSIskOA4AZDOltfmaJ58yDZs5Jta4YQzDvPI
ixYTIt9TlEZdudmD6RVP4zuUd/v2n7CpZRPI3f1GnL+bVlusqx87vO/XW4bXjmh6D0ZslblSY4rj
JeXoxtt196wzlvSTz1MiXvceQSUXeSSC0dn14EMgDhdAO7giULx04o5dCuOUi4Gq3UQiddjJpF5u
gtr+OH+KIPT/vlkRJrPM1aMwfHdyVdaCe3OkB7e7dqBXzHoeSXuQZ+nuWOdd260ApfgBEEi6JH/U
pw0wWHefsSI6VTeSBPpVsDCH3PjwFUO6iGyExzzxxWsttiqtw72Rxe7siTCnjGx5PQO1oR9c9atF
PSUQylWt/yuG81fzbUE3LSgzZlSoYF9ESvrgGQ429Dv3knSWdSPUB6zC3Bk0xGCt0HiQ8Jq86QiH
+LuddKI+KMbZClxG5/GkDeaLdvNVAK4nyEg3I8nHD/r7MPCdTWfkuhRfNokuy6Z6MuIb2E/FM2it
C1P/shLb5k5D41LioraTSTCy+hVoXXN/QrLv6AmZnJ3AEhV32ozKEKC5dBBz+mmfB6w+bxzUkJBo
ojX27JlSTMzo3WaY4B3CSF7CjetPhEoeNZx1LcasrzLwiX4+O2OSSTJ2kitp3hMOpMSmJTGixYmN
CwrptsyY3bCHhB1JJ+SwmBimv4g4eZ+SEq4VeM6dUvFNh6X7N+JKLgjGpR0xmutzuufh9jWKCB9y
YwLS9UGOZlIlUitVzw+np9ZZl3IS4mnVzSNm9n6bVaNGiP6oSbErGA9fva/FAdxjpYtI5mI/whKj
tuBTRoAy/xMTLVSADCNlC0F1C2NnyyPiRsiDkS4eNcL+WCqBRabpTPnzjj9JPTewe3XAXg2LC+tm
aJGmWwjWmBAxY9IJGcpW/YCBir7Q7WeluIqKIDZXXM3822EjbHpkNF7sUotVWPWb+Ghyr7qspif4
W2hTAQEA1WiGqKE16HWf2V3PAcvfJ3Je+ogtk8Zkjx/4PcEgXBJA6N5jRSxzlxiW3kErK4OF3Hvm
LogRRN5+W3sRN+EcrCsMsSA5jvZa3Qm7w58PvTM5aIQcOAHaZzJB/IV21q3/AwVrNT99SYrFiAWh
7O/eizs7KhqsQj4WmwE/a6G1NTpoFb0x49evabn1jWYJ4RIWsJMb3oUpCnh88Qx5Ba7x68eqEIr2
I3aYxTeJvRuR69oLVgOktSn7vniUQ1XG54SOL1jJHIVYhxeoAFY6+pmNyGMVPqjpwr0nspXSOreA
bcc/qGGya5x8G4M1PtLGB8bs1PGaAyvfboMMG8itpLmSmN5Wd6Z8EPirzci6/V3wnWba+xjlfPtS
jSNznUNnn85Wz0ShC65g1q0WxAGhW6a/I5vH++gq1OefFCgjDWOcxhJzZrIFIUatpapOV7PCJv6n
RrxDZ3XwX9LNNQPad0SK8e7uD5sGwsvAvkVoV7Ce29q+/JF8K/cKZI91zSoyG6S7McMDOKdd3eU8
7QxGSbSocvU8G420F+bJh5Df9+7/R0o/TAzFDo6GGbHJQOo7iDlPqhhti1sLWCW94Ulgxzr2lbwX
7dmPmdgg+KUqOwTleIIgCMUNWYqvieCicPaKZi0W1bfqAbzimUxR5p3X1tBjI8w8sETPKQv4Q2a5
eIfRjiSruVBZAqJyXKxxplWdnVvkytuCa4+rYGRg7a1AHuSQBg7MxSlXcOH5sZiGbTGChX0cgsYz
BCR/rTyjpE6S1LdjOumgpqECplI/VhqndXtIpVLG1wQ4f0snk4Yc1MsvuJO2XlL4wqD2a7lkPzma
Jy3gM15Tzru/O562CdgNXacVPf7RTk6GK3f24oE1QTBcaNCOvR97llEPEMcjprFC/R1Yid//7uMv
aYY1yKYL7GA5EyD6sWK2Pca16fVPaBJ3KpZXOthemKWUQJEnqkFv0Wp2UEVEknapq7leC4EQRZ3S
R+EEWmTEAd8d2s5MPETUMs8pqXU0GNNiC0FjSG72m1PbQx+YWBcczLMsVzR6btLeoxZsGwbZZOdT
oLU2ddw3M50NsZBEq+7qhwOpqiwZLETnyIqjD83D/LjSOX0bCcz2e7tTB/POHquAWuyAuu5DmRM6
cuCu6pr8CIokwGa+9mvuF82ksSkIyKLnCy3pkfyTXQSyQHEy73mgSpD/l8H/FJv120A4k+439jkp
T9aN8JDgd/HTUwjSiffAA4TSO05k476Pre+WOeEaojku5KTHlJboYRtcttW4FrDt3+wBqF11+2vG
GjIuvNkSbJH9bjdXWtaFK8nKQOjRdYpVj0ivy3p42Ct7ZS+HVbkR1ev7Std2lYci2qk0/jaQbOJx
dhLqGtXNYEt2ITdBrcuNuscwOcyWqOyjE00sqNL8UEA5MTp/qSgRdF66kwHoXsl5Exo8dmQqnuIv
3YxnYo9UW1+6OAU8Cn8IgUddzj3kwL0PPnqio8Vs9LuahcityMzcd+56yycyms1vz7cCSjLE0uLU
XJfO7+FrHqCgX0cw4o/lvju77IEHK5ht4GjS31uSjVIPJy00TO3ArGfWmAiynNrumNCLcataKEh2
DrTQu1SdYLCrPWIx4W/sUq+OJbEmm8noFt7/PCSCpSad7v1reNJEFmxii7v4rkmb/5X8SuAVnQPJ
IN93n6TsLZydZ8kN9O9bAeyeRrdPtVpNGhv2/sqC9wBBn/nz7Yk3rjRcjRI5p9PRsWYbHj/waSNq
3EU48at695V6KpdEdzjy4gOoNjIzLWMvVaeCvoMcxtx3x3YnLQIAtsUU8oRbwMiWYlLqKj+4kiRb
cQ13+4gx1Es7caeQC0xiMMo1TcZwzPP343x00htRgpGaYyLYDJIm3LspOpntR+MuNlKKOwJrr+4F
YtH9duKhPbbMiJIvOzSC2YF19y94GoR/EPfEE8Rf+NqJm1OyBISPuWPt21If1tF76551WyZDYsQI
pjgYg4Y2sY3o92XjUMALZtwsaHIIUL91aS//YH+fuUHe11Lk9AUINPbWgLWE53ROXZoQsAunfnCz
mjobwQQUP00iDuU64P6aSc/Bg0c+ne6Rdu3/CuzeMpcJPToOqEF+w8DZ/Z1XeGyo4s+dv3quBD7f
g/WbBZ4KGKqudFEtwghz1KEEexqdsEtnUQwTntRPctGyg19FGCQr2kEtYy7tnTlOZg1EXuC5ErVG
nywEXoreJDMj90HuopnN9kJ6vb63dPNNlAmMMM7iGTMewaJvlD5VQAnQ5042A+OlAMSDdTE6ukk8
EyG2R249FXqdvTEH1Ju6JVEWUUUOwT44KagjqFJCsjL0eRdoMEO0c5+U+otC69g907NZyrZMyVru
FE5YoY5iucU4b19G/5rWPxj94lFUXZpo22PMEq9lGVR0EmVW2cEerkzXIs5F1uFsVFdPrKB9SQ1X
NJu6tLZZs6geZRRkqqnGpm07ThUVLQu/fb22n3sUJyCGi49vmKgx7qoVp2AS9NflF/UnwaF/Pkae
uE0G+BHYtuF+XXxnUiCtMTNpWopetlbrngaByVl58OiykuNU2TG0O/J4NnKQAES55Pk9exv1deWq
TEdCx+k79u9iRMR3XgaW97MIt1Ox+SeZaRnx0zC1ivSTj/Neu9n+XNQbF6vVdg0pU3Sm8DZERpUS
EMyczZJn5uogHsajXcc1j0OoEG3B5zdguXYpezfn9pqXiQANy90LidHfi59CIj7/6KiR1t9sDitJ
YPPrlyOfr26ZOFLYiixL+HyBReIcentG9813V34+LrLbKs/fWb1/sTX/ikumYRrMA0Nak1OyBOd+
2jMhiFsDjfZ6w3ilcdA5seEcFquWuWsyZbpo7ADJAW2UiJkHbTNtP0zSwFcwmpofkp0AA5JVT+iQ
/SOxFW/sKwsLYmmUpXLwJ3pepJJWvf9kW//ckwxcGezRG+5+RaAulfDZc65Typh530LoubzgWJHx
6UGWiqltP6I6iJqz9TNxXRBDcGax1msspnuh4sXaHEPifkMw/r8x3NXd/CSdddaWYvdNAQl4r1uc
vVNuQXa4z4nT+5nRpwR4AxDVSRaoCkdpPkNQ/wqqWOwu1ta/IqeWRzTV8xCfgN57q1BuWUVfx0qq
+LykguxOxzHStgbuD8AZzGvQ8e5BHHQ9FWqglBnFW7uVQvZSyaYYQyrPh3E8hog9HiD7m73bA4+7
EmQ/yFs68gKLs0SjEpR8ldqN3z6roft2rfoLU8XmfbJU1gUUD6a07ZjvnVOnpDx6GPCCyYpSZVKI
dRzwJfSMkE4PgmScZMO9NF41R6/c/aeYeH6P2eI2j32Rg7q2uSb5nbr3B3opak1vFSUc0Erxei+G
mKdRIsnnLVCMeG6EyWX2cgPxLkw2zZu1wX9MUoOSdjnC3NLJYgkkd81Q+FT807ZTtQuVoW2CqBxf
MNedN5KI7SphrT6IuJ5o08J31q7P5QF4wwIWPjyuGwfxPhzeI8jVmh7YnynFdg1FmdRlWPkf1bMU
yqONLJpXGGC3pJPD10jwATB/hs25eaPjlXUMaKp/CaT7GOZvTMB1j6c9zpWvij9RDwh+xYIClR8E
GJuC2dCOtzTdObDWYduMfLB8rPk0G4MvA7z21ZMXtiopy+KmaFlkelTJZ4Dm3b3e7FUmFouENeUw
ECfY8pyIFRv9wl6X18R2elkOEcqce/xbh/SqYcdpDbgxiuGGYGgDhqojqE9P4VYo50k6KQC18JMK
WpgEVcoRC81ypkILDtHvwg+NXI6lXz8HV6XptykQ/LKKV/3DLF4eUxNVqgzo4xHaJECHget6WGw2
2wZ/YSmjcjLDO36mZzaogxp5z65BpZy38nbTYWVjxKPMOabdXlpJ1TCPU9giDX4pCTHer9onQuuc
x4y9G6T9SPNWT1UpRAwjFSbCKPvXKKlxCT+0NYtfYRNr/Va7oAmnIEynh36uhUm/3RxXHfia8IJ+
lahIoUPue+k1ou64A4EyHuowW+GORtZWzVycEz/vQzyRAl5zFEq9pgGYOHuClB/JcEVD3PuuGgnh
xc+C/+QN+kSZC62R/CP/RHnxsxEbnxXhq40NpF+obVuEJedrFJA1WM5ZN1ErY3d6p/AsoA8VNV+i
EmDF9BAeqPaxikkBur4x5JoARqUVjvl6XD9/yyaYTr/370rBYjW7xBTtdYNTIkZ2v6F0UIgaJlyM
5AKdeKj/Y7Wyaqhh9IKKYQD4X/rxSBgSyGPIuDK7MN0ueoSHdsK51DoRaYP7VBRh8Q82DL+W1z5p
euPt3I069UTYgKTcOvr/JBaF2N0G7rsru1k1ER1hs1NTj8J4+5EayxTXOg7pQFZJLr0iWF3I690t
7QwkZwORLN2c5mseW6AVEfd7rufunG6P/p1bkSqhoMg5UiGIiuFN39gMwd2YeJld4gmz1dZNdmZB
i5k7cCgXDUkAAciPQm5RACaWWPov7oXBIR110HBkTN3HNPuFc7e4uUZyJQTnkBm0G/X3di7/LYLF
TEH67H3b25f0hX/w8HgF56zErumOalvnN4bgo1l2uf7nWPRdDv9cIgOfxo/dE5XRlffcGmJwWFfF
byVHoSe1lOxQAsK0AxlAtqEH33BFBCu6e0qwM0v2C4n8negrUmy3zxm1eiAhAVoA7CZbdVgqzkpY
+M5bJrO21kV9dqxJ7EuLjBQ2CCt481eCZnA3S0IZZg2cy7p7OD1/t0gvdbODNET09PKxxeYuizqP
df+XVWFy4qR76bk9LCZi0uRCtgFGYVdWNNbB3RbO6fh2xcvp5d2NvAs8Y8kqdAQBmnCtPA1kAS7L
z0qIsmL9WSbl+yoOTO5fcnUbZ9ooLVe6VAwDFszrsGTRl6GBY3FLokTqN/T3qTRiZHcjIou2MCcO
5JzglNSyxwh9e9rFNqwTFF+/0KhW9utu9TD2MW8V+Z2CFS+rlwA77m80cTLDfu+XfPkomI3CW2wq
aNdT6mrmgQvbpKJrFmGVSOecLkYo+8ilHo1TrjkywTc6GwXUDlmq+j7AbA4ilS4uEe8HMCaAWKKq
1bkyk37QOdQaAro+zHzccPc1XTBZ5iotuJsn1vekIMkR98ikreRXi0n2I0SK8o8CQed5Ma9QKdVC
BCgLUvxkfKgdTFR1QJ2J/O0S2sKf1W1UoTc+herW6Dw6dJviryPDgS5cLbE0gbBOwVYY7ukONMp0
rLy1VjnVH1RmZFlQQhZT9Tu/abT9iC33cdsZ1Mj6375nSx5NYbk/VWYq7HTJu60yy1gmK/LrXi9v
15b2KTQXgBuip7crJ9F/xGOJov9lmdm2sBsc6qj6xIoIHqoNl6jsJ7xAVvtghU6PIqdMpw983N9C
6A3t1cWufaLwhACcVXg+/NKGdT75ajS9t4HB56bKjYogQtIwod0TgjPx2mK8SOqN/UZ35B3kqb7D
1vrXayCrdlTeB3KSOREVGEG9wt3KpkI/yd5KTjt7xZnrM+eP7t4EpRxsJTjbr0+nC2wRjkFWBTwr
HDdf8DckncmMd5VERtkzYVzcTXbZKsCidcSf5pCysVK23HhF3gHqahYPNxf3ydrpUj/BDKvAz8sn
75YcyzhDHHAmVO49wP8khy42P0NUs76RRzPNp35fOWJm7s0CPFIt+whVkhF3ELEFb2FhzK14Gwgd
ZYeEyxdLoC/lNW0gcHIGkqWnCZRKm4xjUjbkphAc7kFQouEMz8t5P4Ej2iQ9N+eeQWCqcucyvxHf
sX7F65FCgOsp88dt/5zMzAALruDPFpV4zsGpEasd0N1wOvPHccADIF+ulrFnxoH05CtinM+fwKFH
2WTUdXnBhX08g+TA1iDe2k9k6noamkkN9O42HKza2Iqs78Ye417Q1lBM5KkcJJ3otwXyrKGT5d0F
7EbZ0T14GF9nd6QBSkdf/eXxW1luoAhLC6U5zif4N8wKuZ5waVJZS24uuGUVcPNmIPQ8WQB3WnVH
1J8MxLGZI4C6kyIpqnRNB6owdWiwot/kEbWW6euG4Z+aPLDGaVDCKOufRgJMbygJUHq5LQl8WJnx
y4EwQ2sZZBlxZeFpETLSiTD/GrDAkij55eKG9HBZf9gR8RrKdSbTaiPgyaCsWiPpeWFfgK8BH605
fiPGMstedKg69bHmB5PeY6Kgq45Tr761TZVlvLsoAiOd5EOJQgpNpNtqA5HkWrl7WlkypTwB7g16
KaRb00LqHWGzBlYaUhZiok8L+moTN2r2V51nBRoNdR/J7KfLRYfk+VFd4bT/+edqdilm8B/fKl9P
3D7OBDJMMDaHswB+a84veNwSq6d32yuj8NAXR6PIELlyOAPPFroQW4yHXblEPpalRhA42VhwhU1U
ZSYRHYKiMQHypWoRAF3TFg6eMJyEdcjbtoaAPk1UrwzEPWi/n8kiBzJsmoEUP9Wt84ddDWUmY88q
d7YH5IpJfA2uHYr0D/BzzZyZX1l7LAb1ikMPYh2je7BumxK/mjg3McxbRbU+RJzN4ClIsNyIZsBE
Xh4/NkUCFuH6gHfFB7TkCXD7Hl/pxzdzJvIoyU04jKYPGkyv0jfQGTGVsBcIjB5QaNAw+DoOhwuU
3q+/HsVOLiaNgcsjUzCEu9ESqtXs+dxLbQolsmPBcqhP+eJeo26EnIotGE0jlpR25DqQPGotNeSi
VwYCgxiQ9jF1KY50HziWVq0Wvt1/xmhQYamJh2ybYsDS7mPAzTH1+UYmNlm/S0YUujEZozWPzZvO
R49RoNP/PRRCWKR8dWtGsKi3Jlqut9d4eQztrnvrmmeprkJIZqqVvRySA7cFJ1ETgOr8gGZimUQY
uCzwx0Rifm4js24JqOigRBP9OyDqF7JJyc4DEKgdkOIR1uVzuajupTlcdxuxeYb/qHQcB/w7nj9w
+xrQJtn0RfAisA3F5lunNLsvEAcMEeDRhRJN/3O4PN3MzINVhyegSNbiDsdKg8Pa3Mcih4dzDpFO
TSEkrP+Md+ApX3fw/2NnL5cBzi7CIJ9c19HwV5XW/7cxiiPhH0970Is+zU3dGIaGsFujdvHcXCqM
pczmDKnSZQRRwiG0LFivgyHFt6cgCox9lGBAi9ZXM42zm7tHnf73iJ0l2UZ59PM2m+Gsl2SqTgIQ
e8i5p2nzzh5zUVyiUXVol92cMmzFLKQkxqhMN5VjhVZH0zN+R55JTofYXknnFHRkD+McMUyt7mzW
9IKOkaLrFJIFJ2q77TMYaMTwidarQjAWBfqRKpq66g7QRrjLSAnmQq0nzug9ifRAKD0MxM1wCGTg
6PHhNw86Zu6HN+JrPrL/2Wb5wpySjL72NGhcMzgCVZWqMuRSNP+TBUE1IbqfDdkTT5IH5/29NU74
VCjLEYpSUXpdH7LUP6IOqM5ona/zP1zZ85/2KIbFqX5OMSAeEjQtDz7D7kAf5qRuwhtK9g916RHU
Z5mgCSgTKpQxmGZYmG0ADeku3Bp22CAonBbCTDqmrl5QLVef3Fqfo+9O7x3Zg26PbNU4Ffawf7KH
izHHebcF54T6C8iG+qU6jPi9T0fXPTEt9LfqeEV3Y9A3MG+vWj9dxMVPoeaivSwSHbBSpwM6fDVt
FvHn+RxcflAVMHld4v72L0JjJWXQS+PwCwYCM5HrEkLUUHKGk3CiHplRWSgVI6ApHbg6JHjMAzll
JT8LfdhFpkleAzF4+M8DBGbKBPGb0ClFvS/Ru9jVtkGkrJvXYdbQyRptAhu8S4gC9sluLs3oSWFr
xqSQEIquL/v0/xBEZkIsZe6cDwNs252Q91omy6iL7O+6l/BeTApkOfthRMCQgLxvuk2KiTk40EST
SVYLjqPkiqMqSXcUk1GJH9JnKf5VT/Hbrbits8H00QLX6LQ2z1v4BksvVK7Q9idyd3WuQi1932ut
4vp+YF1r6F2hugjIaBZ+CdxINmqnJ1opCBCJc4lTOcSfiHCViaHI4zRD29zIUmYB+3fqW2qaQby8
SbXTH1RnpTz31BbWeqRAy/FLR2NkWhmedOub2F/ApPN1nW3WTjP77b5bxVLDIaNs0Z7MSYQHA4pN
T94Hr3BJsi7BchaARWTyyXfWts2YhbszR2jdOnewOw4K9hgGftx3bJ5ACf+ZyogO1ZvRQQg4QHfk
McdbwUD97O+qpcp894lF9uA8eCnBclvG9vYaxq6whWCDmOsxkUF9bQJfBZSjZNZ/A6QiLmZLHYuL
E32Ghf7HAAFtIJIs47EZFNRjUSFNh6n4gbgWNkTCnY81BRYM2bE9ZZrfCEoUBrlYHrAeLTOydroC
9V7ObTtpoNjVzKpN/GDir9zmj44dptDq8u5FUxSJTTZdXBOHHmSkYnZ9UenX3zbpTUumwDySbFf0
TzCZxqBfxFS0XB7DepMx6mdziaCg047OCLwI9nWG68x/Vwu7MZx47KAqE7OnHZEqp4IHfFXmyyuV
OmGeD/TLIXskynZor8ay0Bhp/tO6e4xd5uQ7bZkclPLi31g7ajrZHe9bKcTNJR3rQgG2YG+SZ1Lf
LAvCMpU/KqTb95Dt0izWA8xiFhH7hzy1uO59p63YRTAZwoo9VXCUCQkerrsGPPXEnmlDZGNCRA4c
HofZu6z6gt7psbluEG0uRhLUSbBBK37KwtRLkHisIb5si4nX1u16zAPIhaG6rJucgARjjncqlIwZ
LNTStEda9asJFeOeoZMRmz3PiNNMOEgQzdtTqF4gAL+Z6FJXK4Bo9iAdktRHUEvTpRp5OcMm9uOx
XUC3snDrMaL+qp5vq27q7QGz+3sTEEzzd5E5f25TrRtKIpI636eaJU4PCMoWVd8ijCcIy0GEcb4U
FrzNY+BeYVzxavBjO9/jHekfsZnc3t3rT4v68SDrroCqpO/CtSLDh50XpHOvpfppKBtILar2+xfV
JcPrKN+Gx4InR1PswC3N8aIQu5uo6xcBEc9mnpH0YU1mhFk2xdY5ibjoFXrED142u512tl3KrHYC
gTxckzqSfWZGDZ3Yn7z0ZHGfNg0b1jk7Ncq73lehVKt8HsunVNvneO8Zetqc7xr5iiXuJOWIEzyH
HdZ1OUEr3t8k4b8sQV414f/fwyQWa1wh2fZRIR22/O0OGH5UMU+xiV3BbOmJfIwIs39TrnfQvNRk
UcTNj/oI6FGpP97BM35ZhpKaxPcNwl8GzMFGxdsywej02mJhplmB0IvYpSWPjUsz7No98jskcNcS
NHyXkuRld5EyqFwPtmgEY9ZtdHiWnWG5OExtyY89UtNeH2OMLu7iRamugTnM3+eJvmHQTE9SLebj
IOQEJ8luY/cSaB3CqH8yjlRSp0HOS2scYivFnogme2yifmCrvYzuW5s7vUU01ZVlXREOWRno1y4S
BxJ+Ma/MaYWm+DuiFpfKVIcsD0U7D+BQeWN1N9j3eN61mxW7uLCJ4vvxR7XyXuzF1oiEztdO2Kma
r3K7NBMAOxhnb6Pm1PirtB/Svv1G1KdGkPACX7OguDpJqusT0QQVHV+KHrkTBNm8O/bBBooEyGiD
jhXNG+aO9KVyp35c2+6O706rEBGnxFHpBLRwnlYEOUzk1I8sTH8cD5kpO2yGjkX9AWU9GzI3XBXr
xuA0bgoA+MtBNNTDqAWEwleQv3dwlnkrdNMtXJ2UZ3OS6l21ke+T4PLAoDyz4A3m3z6B9FEmEH8/
XqoL6/lCRvpmIwyC5/YgNXna6Dq2yGkavRS4IeYI+7o4eA7WekQbzbrSKjQEyOr2/dWrQz5R4DP4
1oLxjovVCZoRIcThO2QSaYlLx8bJSXyZX4dNsohsb+ooZrt1K8kSMchRBmd/gmGlsrkGOqHZhs+C
bdqdS9Eeo/BjQANXq+P9P4F/7nx+8bXdvdcOFZZbJ4QdqmV8HSiMcquuGcuqes5TNQUdEQPJXjzD
aH1q6glqjiPPCDVlTDwJ71KvvlH9TyGlgk+4fmPxXgWe3kBaFAlqeT6kgaE4Es2EaXL+KU+J0962
znU2yQtNG3cSpxccxiZGEOIFXUQXihfHXS7M8FFAyISgRvlg5pnwcTJGDgX3u87QePcCS9sSBZBh
OIozsSWELgVBXuSKIx++mCxvhtGP0JQZ0/2kP5U6OQJ7QI9W1WuuW3nCrxzInKdbuxrj2qTQUGF0
h8YGJ8hh8AYMbPw3kB68zvPwmmiMAEtierO7YEnu1QA1s8AT21F3vezkMXthAUEcBQiLrNhTBm54
lW+AEtu3jGYTGTDOGvmkQg5lr/Z9oCrT1nlDiZziTGqKk8wmE1pxX3ZvpPl+O41JN2IZFznrHcZw
Sp5CDfwr33Bw0SlcO3xOwQx4gieav4KgBsKHaCm5Y4vabK1zS9pGdOGFC1G/4dGD4i3bywqIYTDD
Cyt9myvnJvi/LE4jYwmCqR0z0d3JJiHxo72FIp1R3uaSopgRLDP5nN+2ze+g1FG9N7rfjigtkJ8R
CE0RqIE4xvCbzxH+6P0DVE0c4WdfIyZyRthW6CpTo38I104pwZ9B/Vq5UMq5w+QO71ZednE1K3S/
5ey7za2OcDnFPkZaQ4v5WmojhTaIQC9/UbmEMwBByPOpkGdXWe4S107QIQ1oKmSJvx+/vR9rGhcj
S4lkZI55R88UJAzea5UdSoad9HViKdV3ydfQVg/CBXJTp6/NSUU7mFgh9rAxfhYMvIKWPbNmBRXS
bXK4RG6+q8s5VcNIbYTsEw2JPbzSKQhoanF1gOsdmR3tDg2LGjDGTVLreAMqS5JLzHWJsxcAof4p
bgzcN4xQc35sXpRBZgs1K9RGpIEg4CE+sKZy9pU9ufciBWNbVUHBwKohTb4KZQBSluc0BO3TvP9n
QqJ+Ix0WVhOlNMmfOvCe3XuSvwSgJlYMgPuCT+/vaW87ypAf1uY4JbHkKbzu/i1gU6KsbXu7WD+W
EuNVe+/APzol/1S8/dZuPJ9rcF+Zhu9fK9KJbdCrvuxVoqkYmihMhZIP6SuG4dhQriSCkh/FVHT3
SkUVhNPBoGJYIfBRmVAUhCGFU3vP7HyEaFNI04/4UP9MCD3Ts9t8dpYOlx6xSyLUXm0PVXeCJ4jz
GUJfVePbmhJdKiVV/cNMpojdtJ0crydkbxKnGmftcEhhS03uEoQ1yhe+XqqDWVThg+guhgInkupL
THct34/aYJkFyOR/sv/eNlmAQcK88MKojGi8WzAQUJHjkaphxSx9aS1M5rstW4AjsZpze2wObGt+
grY3oiNCqcbvQjKukaGxuWDFCUht5nj/FeCjJWa7kbTHCpvD4DP8xvsA9ccUGKexvImnP95jXi/N
D7ysxv+FiLx0VodEfaTU45bp2Bjw6mCh4ziQeLxCHtPzbuMqBY3FRFaVi3d7hOgs4auHsbbdiaUn
TPSbLTmeY/l501Z2XuzjnqDPuWxrjVCHq61HC1Kgnin43paiIW39//+4h6hJ2i2P/3p0IeC/eLlU
KlKaD/uF0N5AbkRQB69e7kzraXNhR6zNmB8rrNHJnAhAUStszFhp7BLPXzzDvhpFa+EYoblGXwjG
WLFvMRNMX8w6AMMD/kgE6k9oUuS+reHEJ22DQXsr4rX7w6g2uG+AQONCoC1eXClFJ+Bv4jQmSqDk
irAoNxjqQZZ/PC3z+36uVqgLeeOik/2Tsk8xmoE5VqhuRHTE2MUQyAYWJ8fSP2HPhes00ixa4H6C
z52nrBsEe8w/HVu6LFylFvMAwcDxZfZfVem0awUVzBsTM6MfQfrHwPAIXu56FpyqQiqvq0QFBliJ
Xx42M5ePEx8A9KuhxDVuf/yoSW31WS55NMYHSBmO1EiqfeEwG0sHLMyCwp+aEJTiPzcyRJIjsoc7
bUYkmUpZ2M6hVwwrrSbDrjT443NJh8FflBcy2thMcIoi48l5Us8qs10ybbpLBAxGD1Pzl3RxVPiL
5fu+Iio066x5YI0PYRK5lj8tyIZyGtUig6K3xauiVypr5wYqh0vCsVjH40ZeuB/OLyqdMt7pd2sw
SItFxruh0yiUdmQiOMmGTa+dXZpITjhlmcha+9PiKdSbpsCTRuPMZnKFr9A6k8fhte7AzRixxHYk
lY0+kVMnTFT5O2irpsz5x9U57gpCT5cap94y4Wgepzuc3JFY44DpG9mMaG463sVVg4ZoJ+FaFqkE
tAzc55GQ2grGq7OJF9Yq83Z+Eq9bnRm69TDUTjl+AJX6E4jzn4HK8PyfaR3O1OTkDxhUFeNkQd3q
v4HCXer/vHZRyYdSRjBNIxzO90Q42hzPZw1h3eW5r+dKWCkLomLpPxQClnQ9sB+aHRcdpMQRzbBJ
/5HLqYw9RrSoRmnE6DHuqlJku2z4qhOfftdX1D1BrT2q2oXjc6mFcY2y5OVXyfMr807nT+jZQvqO
pmCG166Scg9r/GDt0p/nZROR0CKleWyOmXUET/PDjUGPxJdykkuimCCkyVoZBZ4QRSwgSRoyJUQY
X1UOiseEjeDsU4M9XmyJpQtnKPjEKlN0Bicb5RJudL1jPZoukeQVU2D763Q4s6VG4vSDm6OouGoz
vfPwgpAh+PKP1Df+CBYRx8UmGjQpEnWArINJg35FyqSQjpsjL3ZF9T8eiqCDlYEzdohYZkLb2Hqf
K3tqxz2IdxEfP3L8bbMfUFKpgMqazQ08KICwC93KOKHVviP1mEClkZ1deSU+EbAO6V+/cp9OlC9L
PwDxIdRqzjGI6lHUrDqjqRDIxQ3Ej4fj+M1zxeLdKZh7uyVe/6TA9MeZrKMi7Fo6BDPs/0tyjlmg
vLmZicT57QOrCP/u2+ACftPFCMjPZDiYwXPFBJClu207b8gHNMkPniOpqh90XXNZEZX9LG2ibNZ4
vs91IeStk9LTvcin4sZziqvQh8s1EZkILvkrNxrvvJ0W8zNbWL8ko/Qs6nzfgD6HSug3t1pPQ3V5
1qg4iZEV4z6ituq8CvxdObdW+5FMIVgYBBo/zEXsR8u+xXvq7OXE+9O949VnOQv1nb9D3QpHLy1g
FI2LeTbckrecKVNDgi3mHTYn68kLzNWE+BURcqXuhY4jBhspTmYiWBatK8X9KkGUUl1uAbmotcW/
4apdj5nkjJ1lRA+qG1k8cD5IzxKSt3CBzbiZcvH1mvOmclNqVIW/J2zYkaLrCgSeGa1yHuQpZKjA
itz+7SSwCVX3izNt2cuy4hgf+KhOd5bxvLSKoXqcQgocTshsiU1JVed2Ij/LQ62rIbVWiybeG9aR
JNpT5cV2w/86EAiMehr0YViqlG/CH9zFCW/p78TEpq2VZyFxmwOEdi4rXjxuPcbv9WaAkXaxUvtv
TELakh2O/UVMuvbyTs6KB+DHUBL/fJ7VuqrzRF/QBpxCkDJmq13uQVvyEL+6YYN93vfbgTJ4zbM+
NJ3CoFdRK1JyxyxJLOh4ZJ0zpFKVEaB2tovwUD+wf8ZsVUJKG1xFW8sGeI2TfcqZIYOKU9p0Egl9
gfshVs3hg3prY9jaBQ7cZEbRucjylOizW66aHVR6QInHD8QR7Ohc/8K52a5AWbLmIm0S0lxto+r7
+SKz12j0+8+78abbHCWFt46kaxzgx28gv5H+46GGrZcJXQ+Z4f98EZ1Qj1W3qZk/jw9K5L56f262
i7y2mUqDvyigOdymfTSBLdxAXbZ0x+JMVyJr7/gVvN9xEG3kAY1pMglfZhEFUcr8g+sretDldQDE
2+Gl6mF1ohyooKK5R8NkCGVw51GXI53aSrKmfVyieVDsy5qGUJo1vv0KF4wuLICJD9ktI9NXaleb
qx9GcyZCvx9Jay64/7WZoPp1efvAlF65qUCgXvH9jR8vEDMQBCIiO5Xi/sjL1G/2zaOoJHq01LxG
JbZ5LHQe13VCPoAh4WytR3tcriqrzAn7l0Rbt+58lx61EOzE2+T5oiOPCcePWSeoCliSn/9PKGOO
8jM9W0aYMmUqQf1K6nvEPg6ZPomUBZ81PKTUkUFrTJRZsIuTp1O97x+yr+sbRIU+u/RcaxYMyrQl
O9uf7nCdBZAjV+jetaKZPGt4PTfqmhGhGlFpk6/KUAFiE0cX5ic9M1Xzv7AwZWrNO6khrAAkDlhJ
oTpygbLACab7Ctrto8EV/XL34jsCXJtEn9YLMid55klFykE/jD2HbpKXJ8VZ4uwsai3JYmN6yuSE
bKlJ8Ly+4LuwM7Y+U0y3brRDKKhEZNTu/b1CwrVU344kzdDzKk71D0vjv7UZeAmKhNn4Abu+EO0F
s0jJVSXyn370LyfHF1Aqrc7gqHKPHLy79yU7cXEv5CQvk3j7PckVRwgomAFG/2DcxPDWTaaqOPrh
LnUs423IYrN2YSb+U/r7aPRguJn598mrCrPfh8bRkVMFt2Ra03e5tjUgao8kmIKxsBGVJ2afLHxJ
FXw6pQ5vPQwdEDdckQKVkhrmVJIQWXejoP/Tlyf38B9dP06dReYvYcKpb3eFzx1+ThDCIYNuq1VS
5inuhOEa5kEKGOM0B1AB6wrSUl7LdcpPZL9RbDosO39pA6WPXmURxy3J2XnIoPNiYSfes3XsZGlF
yHkkAAzUx/uxs50phf6ZA0Jlcef/0FsOb6bvRNuZRxVhIzI9/IdaeFQhODypaRVZZ6rmLAFo+iz5
HIxYLtrEI0n8tvl+Dk7fzwOKhUJAz+nB9ORVG2HCTAmR8m/9EgD80lJss37d+cPcKK2pSd1gUk44
LKC/rgPghx9ESxfHih7bJZUp2/hIhIJ+/kTrJiRAs4HFm4bZLXLhsbS0E9wWcW+wmE0mjPXkusOu
doReDnc8tU3UsLs55MNoOlYwnp0iimh0ZCIOHcZsUg5HGOfvxNQyxOrO2+ZlLUQk6q7cPYQxSvX4
yJxKTGj46le33GR+fBZLgAHCuwmcc9l4YoPTRE6U3E0xVvbmPLeLtNH6fj516Xgs0BqAaC0+VHCn
aY7BVBP8prYXV6WZ1doThLRkEkXVZ/JK7IkdU4iBnzDCJvMuszzqggYxj0Ke4G913lfc72lUSKHx
W9dzHgNKb8laOXJrowIKmyPZuqis5yCFgdg2towNJN7VjEBKPJVrRA4jZbi7fVI20Vry+WET8xPj
GWqSl/R83V4GeYGoE3V8NILTn0c5QgrP3C4bUxDF9eL/hOcKbA6WlxO4kVhxP40hXQL0lf/nQnAQ
5TOBkEQq8wseSDMHG4ncBSdt3oXEAMUZq+NFcyzZFSSneqYSHGQXaTi2GJYPcZ6ewA+fJYrnmiLh
tQnVu/6zvzbY7cmmq1zp+nsVNhnOIsU2E5DPRLKOchx6Y2zwLfkXUQ2exTZC3Yfie0vzUq3xuPV8
1x/xPLkvBx7sRU724if0tb4UkSV0zqtMpX9e4cFGmWqLT+PShEfSSEA1OEMmevBFaB/t0XoZMlU+
zQAcoxe0z/xs+MrRRoYpPm19FJ6BmTZ3x394g/o9xpA9hlCGktgaBRVPG/5vBG78cdKsW173RsJ9
eqzsKBBNQv2HBRsKX5lOwyPCbw0bcRZAE9GItnQIuZ2Jcj03zRHl7OXLQ0u2MmOcVWNyLb0I5DgD
U8DzFH4uXjxxGVL7B8fnhXLYHVZklbObstHPz/6vkisk21rCc77XbKktRxiuLY9CQKaPO5RcuXx6
+62j2MQWkOWoRRyx3PNx9M86KKCpxhfJKSc33zCYaazeKS5EHRbTG4SaJSnz9RIKzGOEMIGpzBvw
ZaKJLDQdLMRbdfJtEm8g8XrAj13HrcPCP/YWd+IyB+WRCarBTfbueMt50RwTKlY6uU5oU0xD4MHP
DIKRNcycO5Y+IiN7q2LRdai+O7qMpgFpS0p37/D0T5dxJoWk59DnUCEE83xRw4cR3hvX2mp07bVi
732KPm8FhGWT4xSNGRz6/nPn05iESkk3zfHF7+8U6aXyicB3H4GRZ03usgiJ8+9/Zx7I8cbB6t03
rK75kuFam/l589AJmipJp4Ur97YxluJWIgKgLyHUIbxrIkxP4mYVrXHtzRHJ02rjsvNGAyZLvA1U
sZ5Gkf6zn395VyNxEDFxoUT/Ysc6c0hDoFQ9gp2H1oBov0VB+vcYsM2Gfgz2rj6p8c3Qu/Ey7mju
wnp79bGcagt98OxSSgIcvtmQVUSM7BId2RgErFXI89Tob1A9y3NkoILvUjxAZN8+wam4x3PHE0ly
WxmaDy1SIDUDZ6VPgwvHEzhWwaUbyBagamtwQb/pjwQpZI2zaDALtBVrbnMUzUA/ICl37tjF3FFM
A1AqRILVAhpK1+g9NrVwZ/zjJv7DP+gc/wXZ7u+UDIv7LikRGtLSdBnvRXBR4GSqtB2F5ew2FwPN
jDLUv+9OA4TyRjRa9x+BWVo44Hvd41AHANc3Noo7tGTMun30gowpwN8hG87jpDSvxcAkeLvJc/5A
OIM8GAmuDSl1BAL7c+0WkYhofpd6I0LgBeCfiwPRaweHw0mhuc7b23ZSp2i1QV4CKNQZ+F53NWob
f64f75iIKu9u0iBiQnHDcYP9a4MBHLutpcCnAt8TUFRTK0XG1UXAiXkUufLkZpaho0OG9JMbKIJ8
SgjxxlMowk/7ZC6R1gY42zLfUO4Ks/Au1AsECAqoKlzLOO8nUcfklAcUnhvRsaAvoPNTX7IClyf1
9QHg8NCQZ6oB4ZpQOxi4i36EkqxKswlBU4nkwhlUnDPqYSzfq2IC9uV2iVpUiVIg/g1jw6X9Es3g
wyC3Aqc0yn2KLDK0n9WtNEvs5rLf/EuyLH0RJjjOrVgtwVnlx0dlvZOZQZXyReNCiJILlj1FsDs9
RXbzIidHtpsySD6iWAZir8ibmL2Bi1uBp4sm0qe5r0xipqv/yvglYbyaCRoEYuYxO0ae7bapqjgK
VgUjp9a61AEuGFNA2hf3bTZ7SkTawP+R9KXghPkVNHVvr3JE1Rjjig5MXd1NPFhkjjmyTuaKbZiP
vNe+rbQex+fvA4jqxZmYrvd42IvGJVWIq5z40BZoSBvxkVljxfiPNCO2OMSqepTOWX6P00sBWImj
AMR7Lkk4kwkEYLMbY79yzt8xguR7+baX94+lNqKFtKxCYcC0Q7gdaeVbqzXKeBOE47sA58BAbzqU
dbDp3U2tv802wcoHx8uH/Yovp8MMOQ3jSsMhUU972K+0LGJuCMChI0xOjz/NkwDoSugr7eTPluUR
LFBMGpBh2RLS+NprT1RE3W7/UciSbxDuWtSq/Ix776sYvcK/cSbxHmysJ/mM+fweVyzcxG6FD9TA
KAH7IJQuS0yA2V0ntbZFWYy3sRcsd2Pn5wu9D1838RpHlLovVY7zXrg15Y6BcsLpCea5ht6XfArs
fHQUGt5oQ1I1wws+EbiozIiVd9lDEuspwKbs6Pq7RCFLIcpqTtLCerov26Vi4Ajia7TMjhIM10Kc
oXsPriQy/u3kgGI8P7TA6Lp7vtAViqGBd5BJJNOJ17FXmVYJwNB4j200qCXU2dDWOw+ej8CgjzgF
x9VclmwvLxExBBYtiglwnLRAKX3MilPzk+RsDFxdsLj84bjRzYULiMLiZgIRie7TMe0Oxuaa/e5n
B9FWopEwkiSMyTd2YnoT3T2a6ufuemWLev06VaXLEm31pATE4hD756+e2MkDoVwppNN2XmiTqYWV
Ur85vQuH2yCWVM4Ef/FrJxdGvMFWyCWQeEFjOvy1LeZPLO48t76SA8svaPqwih6BsErTFQmHnShZ
RlQJvxs6GSyb7UcyXPlEMtf38dgtK67+gyCF04NXp+vCO/A2n/mZcTW5x/YyZCcU3xdR8E2z2Myc
CcYcpwj8G2sCITpIz9qXE5D8CJ3mvq5QLCGrmDqCDtF8wlg/LGUVzX1qOvlD0ke9gUQgD08eitaX
9/AcSBuJLehhZcHdc11K5GVg24ozGd+TPuWSFa1LFaFlGNR46oqSjbV4TFWbnXVx+zFIrOLiSztC
Msy+Qn4P9HG5jKCDS0yD+NeZ2f2SRXRppvu7HWCyTOc00MVsIGjEhgitcMfnvEWx1lCmYIFMLWOS
JDA4IY0mO8CUjRYcfOxU3cqWkwpJg3wzhms3Fw611A2XPJv8fIiNUDFH23/+7fJ5DJVxJr+vYH0D
HxaVjDVgTG5BjQ9leZnlnfWvTBP94zML8ywZ42itenoiz34EsNNuUH1mXGZALqhJKN5JrT/MGgyH
LWRBDcIOl+/BUIGIn836N11reeC82muRexYPSxUrF18WsUJiiazgwzwbXQhL/ehkEvXHc7nFbkJv
BbyVAtvzGsikX+ex7IX0BxflN8x8aLuO0ItJ+tTpOghqUebVdXvGf04aj+QUHnhCCt6PusfVRXZ7
mtNxEVnYyxADzZfgutjFU1CEUqa/zZjR4OkT9vdDacUzNDCMtbIUUHBxMvzYQUYSdjvLVCnqKZg5
zVJk4xzcqEKtfsvZpHTWWQ8hq9J7ea8tDZYct4TG9BKIgNir2RktTYDpj9D2TYsPyMIVdo2rM276
+NDmsHzpKW1Jta6L9H+zfqU9sjbbVdpQytOGIpvev3Hc7JPqrugxvaX/hVhlaj9iM5B0NXxxRO73
IWomETMeNV49HOb6GCH8/Sg6X+xFE+D+WlhR1m8GrlwxgQie++rKhPJ9GY11gF7L/TITx1PQFXx/
lgZbAfJNszq24Mrr9zscuMR1sJj8jSqImpmr8OgGZq7CIvZYB8EZa07SaxrSPccbWjItVRPNmG3X
W2DvCVq5WP6FLC23+SELxUhs/tDz35yk6o0nkdOImFXrjQwNoknn8l5C47PV5zEQ6O/khwMjKJua
FViWg27lWu19Q3X3kyP9DOZqoftmeb2BazoUseX1GcAftKd4fYzSna4u02Az6Jyd0knZ6nlP4N6p
5CQ2yQLfn37HC8L3+fooiHgxX4TCWvSvj/kMTh720pKsNWY9jWZwiqqvTkYmUJ9sX7/4I/b6O0Tn
PsZmgU9Ojdw0qyKJmeQtvg7f9Aoeb5tgqSCx+mdfcfVBTzKPELxTYk8cjCQe6stS27M5xLuCZmII
LVsQVsMcPp9921mKsFIrGZLFdWsAv7oqlYadRst99L8J75ayY44nM5lwJKn9hwao5dS6fmYy45fz
DU5CSnqV8KN5Ntjgh9T21vVLblWyIQS2/Si/ID/bKnTpfWAVc6lzs2hVhRSDx53NGju9tKzK0aSS
tgRn1Fhoi1PhtgzwtVg8YlTakMGmMDqWZJp/ugt04t5eVUAg0DQtwxh6XWRXkfsENy6uXD+3/itK
o74LNkZ2lyV/HovHeVZfJHaCnBq9smgUs2ro/44QxeJYG/T0xXmS/tHAgcqiJbTKUx2Z52Io+wXJ
tf4H72dokhCq92NkSZPtngrlft7Hfk41bbBkUjkifrbBSHloteoAAV5oaHK520v6eRaL/VEX6NZf
qZPmKRR9D3a5YaeQFAWu3Ap//Ga9D6v7h/TMUzt5Vd4xi1ckRJ67maNp+u/jrishP0q/hHxVvlf0
nNMt6qEfWAwYvS6aSKelb53kC20AM2PUu4s9urvbXAj/4m4AkienYXIHWF4YhZ37O7hLeYX+cZkR
XgUMZ5QbFufnLf+3iwSOGAmXOr1MBPEBv5UwlEsq83TTvJH5RKwyHVhKRsQ+sZoJLwwY1QbyB+Gq
R9pLp3LnbASrWHEuYQN8fmQHc1wVISv8zfyrvUcRMgRyJGCbLVVzrchvpjR6tc14sKMLm208M3G7
WlBO+uCcbN8+0d90c1FDdwT37kW1nzNRSExjXjz/EvHNvodpiEeVT2GtOQlj1eu7qVVACsOu+EqZ
rKwlK7dT6R1ImJJRiGces7Fpn60M4tf64At+9Zhf1uxJNpcnqsMgjyJBxhWDhE3MdusZQTbukCe9
exndgycyqdz9A62zg7tl36JSUkCDmNxBuZgz5QROhNHnwb8wHt6b/4cXEaK02D8MdJMeOpw+OVgQ
+QU2WpWqkeUuzr2w7oXsbbkHkhnDW6p/d9SS0/8JiAl1equA5Qa0aBLFb3KkvYo+03YveXYOmfU0
y9Awp+bwF8WeiVG1PTZxdqTKv9VSvCppQdS6u36SqXva0PV740eeAA3EgN9cSbsXK/jifJprImGW
L86WFg46K+EH0lB5LCpW8TO9aiztItSh80eb+piVeKZlLBmacqj18YdXYYU5QGrK6+wA4R63zxCf
cLMXMNd0aA90Kb1rYWUhCONEjoJD5i7ZtXDh/IlVlojHQ/F54pgxiUzGrVaskYotU/q6I7eqinHx
Fy9swJd/oun85i/mmOU3XRqPGtBMHL7E+K9XQadU5ff2wwwhh+Aj2Dh6XNOLooXiL+NxD/7CBj6J
JnZB8/gyxoYTZymmAEGSwpeRhiWgLLemKX640Fb3OFD9Sy3qCsSNhcZNxHzYGPrkDuB2fCp3I4Hx
9BvtvyhxWIQeNRWxHGsXWefvdb34c3n/OT/LC05koXd2YXpTfvFOlASuZBi9+4xOCt+rvy/kdos4
qUd8KPnpBsyQq0osx+U4VwGUPOZNOWEQOL2o9MN/h16sg3uVoEW9+Iygm7PHopBzt5TWlVR0OlGH
ujeXub77q8i4yAeiUqoDoitWCvRqRyiTzYqywv8RUZcIhTq+DcQuPUTKI4gkU4TZNldtC0SfCUMY
i0QzX1mxR1mDihzLnsoasPJU4wnr07eNitD+UJqOWK5MzzzRm7ZMu+ZZfAFHR/7SBTZ8xwn7L3oa
+i1ash3XPBiGybs8cfvqips8L/mCTpj2Jc8uwca4MEKQcscSsUBCzUwg/byjquNoGPxW38fp1IWh
rWbyKtrMlfDpz/bFZz+KwCV44PLbcQtpGDmF63V6AHz+0Wvc+wiPj1mYEPSqMjSFc9t/UGy97Acs
ACcrGw4mz7dBnnPe8J6A93Lwowsk2/4XMYY6vJ98dmA7Odyp6lpd8p1gWtSsqw8f1ROuFnGKAwqj
FOgSEPp5zcb19tCYZ92qIzVPTeG0B/Nlp1DggafWzJuUowvWovrZ4gurxq80ids9JTRif734lNsH
SysUYO9/ww2Tyd4KDWq8M5MyBdxfP5JPEUeockyxeOCEioH5RMYTlxhEB4zhCgosg0ohgB1I4/1z
F4ewgOkXs02K7uy1fW2E4B8Qkrwi8hR8LEtOQkOfhqQiKmL56bAu/ba/0gMcpwe2Vw4xd/Vd++qq
NphXh/uYVmnndWm0vDaM05zwbfcCBvZl7atMmcO1ePALtREKT8nNos944TEf2jfmRiDGnbwG9Ngo
DZpkgZXQ04yVVaOQyRHRn+8fV8btfTGBvBdCVR7AkuXM6sYv4G1WnZ525k+P7CWWHG6/y+g+QXzq
Omhd53WeOL8fHWwGoVZv8T84b2tl5czzbbQHcV7ATFGb5Ig+hTbQQ51N9ipe6uHi4RLLssxYC4Ra
ZX4HyqiGrKBOyAmG4j5ZfFLoTm4FdEZg7nlAodGlZqn2gbkXZvhonc4rAZ2OGClGAcY7jsADao58
/UWvD0JDI0zFm7uq8lrjza8SjT53O53u9Y9Ghup5HzYh8jrhkvBN1lhurfGwxnSz7mixxNhB/7mT
pOm/be0gnXqJjv1XLGbipoypKLkny1LoTvs2DeYPKR2YlkfJRst+lYHrf8KPCgGsD0TzZOEcWHnN
k4oex+dPicm4Sww3D5Y4IPidulxW+nGxjrl3oOIhV3Xvdn+p+3KOnjUSI3eAJDe7NxqWT+25xc/S
O9JESM9lJ+HfPmLQdoFKPjhnAo3Etg4DjmzPlV67pRUyYe1w3QJeGvWOBihT7+NJSc81RjIBujgQ
1J27kd6LA9JHGC6nfX7TWs721M/Hyu47Lz6lxayN7iRhk5Whzor0DTr0iEo4QvG3lefRfYGi3pwh
uJa4+Tai7Id6iaV3xtztmUV7313AvRWGrev1vUEykKieu9PM4LdrXCfilKU2DrzCEmZYIQtVAwgY
J/Nct58oeKRYkkOqDX2dajLEHWbZIXf22xkCK+03DK1JolrwmqHv0IO1U2S80KLxobmRnrXtbp8j
ew7Q6Jx8qTDJL31dczI4U/qblgJ3VokJG/QcM57RjtnjzfX74v9BbN/YpL2sOj9jOxyLqEFfZChy
BasVIMCHZTVRjeUVO5JqWKYSFlGmt1tQq99ve8e1vP+Ig1h7VX5sxMHPlriiajDFFgphTxEi9iul
Gtpk66MAUtMIbqmMXQk3Y+TQcFxMlCv1Xa2rKsgythtfieqoWvjhRgMiRFqaYAeWCPHUV8mPNHuG
1cwlLfQAiEkxkDy7vZ+jHoRzAm/pnjbmvSV0hS3qiF/E19dPf5VJ6tJDOaFVBv1wqx0kHymD0rLG
S1F3gdJVucTapqq75x2v/R8mgaK89mq0+4PgyQqIibnzizVIKSHC6Hsa1VPQVELTIAV66bx8HQu4
sLYMBVSdpScNeCDqB6wmszD+7JyHo83/6jOwjxpQNMFqYnLUY87w4vT1XazxHmtWu5XYHzWMfAS7
KXb74BSqsYoekv6sYfcE4DbPtMS8MkmQNGhqHeye9/obpeTh84ESOet14JDrB3LX0F3HunrV5ujK
28CZercLzWsQIRsBJU8ekoxP3DxF5pkdDMNEgd7ghIUs29JPf6eT2XrcwTlbWbEd6QdqbUvTpFUn
M7IePTllkuaTUp7sz2gY91EkVvUcXcXmbTYpJGL1zq1vrt8ciBdFQYc/WpvUF7y2Y5/aP4AZIO6B
ZNyTVg2Rz8T4F3SjSg0Qhz9LvLU5Kx77Wl4QFs/yDkMnndb0gT/eODZJIN+tz+4mvBURd0zBVXdJ
LAunJOYc/vxG332UI+E2a8wkMa4Q5c4C53D+sqRDmmEM/065DYC6Dgl1eLG3yzz/fRLorIhvduco
j65am3J9LQ9mmuQbupJ4oxc8LCGSCpiGyXJwnnzrRl71mcY0hox6w338m8O6I76z8toXhhVEnOvE
OpAn24oKUHrhPcVhwsy9fHdds8sXRqgWs852hEi1mE3HeuMITMA5/Vy77uqGoLl/dC0QmI/sJjsA
lNjhKAhXlWGXjHy3bmBWplFH+eqjonBQm1fT1r+bHJchgP3bvudmw9v3m92HdmqOez29QhZy2X5H
paey05r23AyQGqpSnMHYCCgwKV4QsIvqoGaS/n4u/LwoFRU9um2qGs8ewjQZ0UFNF7brWJ5SNgUN
6txVy3E9nsUOBjnSD2jd/wCpVnafzpCHNsQ1oqIl95i6VYM6PKhOkh/rZRNtMdBq4hIiQVZDmhWF
sqVavY3f5yX+t3JN5KgHJuHm2U2qWmBros9kGPmW2DaVvuqpBI6PMEjWYSCCaY0p26m7OGuK1NSz
vjlL7J4nlEWuOt+2fTkyisAVWIDcdz5p7tCr73zaHSoDT6broMZG9wMMVzojJPEPhatSqxRnNr6T
UgJDgw8stlK1zncQTM+/RpvJUfTRicFg7GvcYD4scqOGFPAHRFZIxhzufoEfVmlO/FshO8Qt9EOX
e8clfrcimSUZuh9ldWVM7K57br+ionbMCBG+tde+Mb+xhDDeRUYdy6FSP0rKHc4BlYHz0mRjjLBX
uZVfQmfIoK7pvzm5ktTpCFd7KPJu0LVBUCznwJ2dbMenwfxBko1hYy8ocoZKBhK1yGOTBuI60Sm7
G2VsPhkuPDy+PJl0EfK4mvdKWhERDwsTRHqmFzZ/gSqfrHpRQkHIiElTETrbLnSYtGL7qRzKzqMu
MFlRVeFSA6nSNhW5Z/WMGcakwXR/kEtTaC8BKLYFIaqmOR7NXYTd6Xv1VGpbB4PhwptYhb1lbkyQ
+dCRqqZIJUB7wbInE0MMHGwFYtEGi7oOwZEOOKR6b8Njj5VjZXB05aeMo+DaA3P0zUhMdhr3Cmuu
iEf0yS71DKWJJV+X0ooJiaf1UBLf5FFtY8bRbZMT7yCN482gGEsDTwr5SHFY84Z0g9DypqguUpJ1
7ka9F5N1yeeEeGDxPlvKwFpQQM5yUWC5RvaVKO0TWwspYBIYfZWFK+Sty6DH3RRWgOVFx6KMZChE
wCB8yEhfoa1xLt+6IherwYc0/p/URT/ie9EBQw1W7YXYhLJY/31Kx24k87aXKDub1jJeDQOAt2Im
KWVL3hCv2G0TSVNhU4m1g0cTFDtRTkTZcHGWwmjN3gc52keVvDl/IYOjvObCZlwmgyEDvEgIS9bL
8ptaH/o0c2zLi/kY4zhslUv/k/Nk+wo70I0O8mwx55c8UdRCVBJ1xEXDqXzahrnaoGTaiXbx+nyY
Q0ruRl1rsv9fm5VgvFiMz+Lt8LaleQKk+54gAlccLPL0teeBioSRTmEgzLaDWBRq6Bi/PIDrXe+i
ToVw43nK4skDmEM5OhyndzZOnz4791a90XNsuJ8XfPg4rUOYLiHcpKPUX8pJ8r3rBeID6AcJhIIZ
u0liOatUMG5TVstGllJDe6NAhsii4RXnnKu5jzcIRZ040f4rdHvWK4k4/YgrLGoKD6T3zPEY1g7d
2KIgm6tYcTEXcTzE+FNgvIJJ3l+iTdeJwrUSj+lDtmL3+wvv7REq6DiKv9qYjc0k9YmsZ/sWvsx3
6SUEjjYUCV9SOrvoz8m2AFk0Yp8kxqXPNmPTPO59ocTQjLS+OQXaTUTpBnfSqtX4W5vKTdQ02jQt
Zvszq0eU1hV8309sckHTo9aM0xVm0BUC91BRVjihgK5RN4ayBhFPaCUS7TPR/9dDUAEi6X/Iikbu
o264fYecDsTN3F2dSI9k/2q7oVpIunu7oBFlIoS20ZOzJoLI/Fmmc3+Dt4pTu5oP3MqMO5zVQclJ
khv47B4fFZX83CVLsXRyxP6KSl0tk5rSBI2/4nopsQtOqmHqLVDS3xogLTitdWnCAYFDl1eHsbSF
dEBXGnndtZ3dY6r9KPCjzZnHwtx1t3/0pfn4AGx8mbdkHIbMpT3x7dQ65bVqlpARhjPbDrThO8Kr
XfvHFLIAh950WyQSRjulV0Q+vDst1aEs2btw5NakgyzRKeLfvkPK6EjruNMdBriOpTmy9ngVkrw4
aqkDNhHH5u2j1F6h0UOahIUIv3Sq3HLhcvGei6b2j859cyZDfTMAF3uQve8+R4LhHirCNVvrHQdg
QA0JOB60rFX0zsuamoWb/e4QDN/uLj16ftdVGnfezyUns7Jg3UB5Ik/D1K91lFjTWvpTbHpWweY0
Y+20Sm/wmt6p5rOetxU0oCJ7J6dngUOvwZXxsDwb6g/cq/qYthvi0r7yztO2h8SpGhYHwAKW5unO
8lYbW6mC+71dQ+ejuaalgxSWi5sNG0HVJ9fxlq8meaVBOYM4kLhMZSyrxHIKWsqeHJu/ytuKDR9H
hJRsFKMkGAUo9IQnye+6Sn4YHX31Q7tDkRaqym1xIlDN14Ml1PILY1Zc0zpz5MNZDGfT4ga2ae3v
xXxfolAWaB8+5BKSNS2pjTyK+I240B/K5dxOO1TQdU934cewP0Y/npBvkNm23jC8f9pViOxsGl/D
2AK5mP5IZYhB8qKUHm8izwFOpja/acBM+igyw5W5sReq7GmUuA24Ltw2PS5AAnOGy+Qud34Cp8f1
preVSXe2hJHYbUlx8m1JW3jpJo6kB7P16tbagjXzEI43jerWHhP49fveXy90G77v4gkKGsm464EZ
7HQQoTkead8u97Oe1BjpPYX06sZhuL+3hQ1yHbi6W8wACQUFgaSdjkcODrU2hYA2I1UId1tnmwZe
2qNf3rRxPY7mZDmfDmQmdmQrRLuEsv1YlKoR0+snMLlGVhH4PU/GjbQ/mKtyDTCGlH8cM9KeAxxH
FGgKDoSWHIkAOf6btW7wTD74ztdBVelkQ45N5iF9k4j+l0GKMGBaDoiuP4WaWibS4jlM/EC5HXPJ
axV7cKTQukR/F+me1ly0npyLnSdXxpBjeCRZn3W42m+62XwsPYLCL1t5o8kz9n3G/fnmsp0C47s6
5CXJVUHDryMwHCBxbj6iMrgfjrdk85xcb/IimrtQJ+PgwcKH7qVh60vM9OVaIdjeDq5sjaf5KCgj
MJPFham+FHot3xb/i2L+rOu8M5+YperDFaB1iCVS39visXYCQZFYpDgq4It0DRWcLXP4odu4Caw2
+wb0MY5id+04Wtm3rUwzT5y8UH4NmlADqcl6byB1a+zKd9+HlgmY6vhqmpPi6/qm8KG3yIFxvM0p
LSfz1vP//dNuBKIWPx4OJ2+eb44wLmYEf/f6bUfURyB0AhuZEzud62Fdv01eDoc3rAXGcF/9+s68
HeJzMxy7vrSnR/X/sxCV4uIm6isRsL25MvS7A08hCNQn44zfgepE60pFPKYzOlq35iXYhpHdj54L
eL4TssBcMSpwMfN35G3SMRa24i4qxlaFcTiezXoYak37LXy2GB8Kd6bU+e8+Vu7TSEPz67f8FDNp
9q8SbOgHz7+bIuAC4nqh/43WslcvWvD7jp3sY0by+owxHuvhXK1UwKXaZEnX5N1A1pi1bP2NGYAN
XzqDtFTN4dthGBGfXAxs1rxPuNJ2SwYfVV/atJPTKJYIB0djY3fzVc5DP5dpFrwthnXUkEjUMGgR
umf71K8+TDuFDVZIiIi6l4/vHtZO3v208oZWdtHhQUiLMQ45kfJtHlUbhIDZYE+r+2m79GqgtBlp
aTddLBVgJOKUFI7Udto38aU66gtxXzKsVFfSTlG7m+aXqkLqXsxbKABsRzSft4ms6tVIQutekqpd
uoNczJl0vcZHdE6PgK/wIPvc0Mjy19u7g6VGHsFzQ6t7hu3+4EP0x7fDHq3x/4a2CmijNivHqqis
AL/FYienuGyPxoOjktN7EwbxeRsE6yU40ZYB9bAmcUF+geIHwgEM+TVDe7sAAmhb5iEuzrSPSx/a
Ktm77HwutLQ3ECOYYslTWX0eLFje0e2tUfJNbulRUSM1GOPzvTcf/HfQXpWsQYidmymHYzMi8HDb
lb/zzc3wYhDJvY70hEShd0W3gIqAMrl9wbIoRcO2JzuIbmZSIGkWIQ0RVWZ6RmvKqd1vv4jCg5ec
B1wffc5hmqO92xL8E/TL11ejTFEv8x83L7PjjXxPGr19y3fdqbnTO8r2YQAPc3Yg+R/S3aPl8FyC
XfaaxJUMDXSCDi122nONwZavcWpejTbiKZF1avWhQCJ4/sd/0cL61vJvaYTbG2Aqr10IZSwDLCT/
72yRcOy3GQJZ9baS4aiGD34nsMCB+agnNEhCVEO65+xw3EBgfXsXOQwWgc/Uhm//r/UHrfOJtIFi
nLlONQ37mEeqd+p+NiRZIDoqoaUDShoEhlkfwoZELqwEOLtRerx7Q4YHSMl8V/vfkl5Z8Vtj7Fbj
xt329qshzXu+JFa5Si4PqqGrd0AJo6JmPoiMZKjjB7fgkr9jfhVD+9RTk2l1uTlpnXshmDWjbTXJ
QwHae+XwIbWJG1MFalHX4nfCmg3c86NW6PsRHosONUSpOyZu7KybCqGAHZHpHW1VNjyk1TRpvh6o
5Od2/JnGTRLRrNfUmdDnvtxZ7g+ouVFLg+k3Wez3++qiohwjiADpe90vi9b7GMPhhWw83iLEYUKX
vK5qJiwqV76F5C4b5/lQm/1FkVugRiedkfoRw38uTs5zj1W14uiIi/At4GjmdBhEvHu6oGSATmji
UlFS+1GXYWOphG2Z4aaLJ1M2ZqTbTqi4w+CNb+17ECBKzxzS71o0fkiM7DznD9oSUksvaTYEgdqF
1jB5XedkpKI4U3F5g2xwymPz7slmMiCejbTujrrCjg1bbm6Rct+WI1NTnBRANMFF5212TVsRcV7c
nNuMqGPVupmZjyF6D0/KH836rWTNN1uRhlh9GP1THt/zdUP1/RI042sYhTWmIwvESLoNI+qUSwYC
MMV52Zfw1/CraIxc8rRpZUEx2EHPk1Z8Wo7IyNDWGfBv3qI6oEHucbf6TCG6vXEGzzaVaBMPFKht
o00+Apd5bLNvw8sYPjZZHe2vy2DjHiJL1WnW7VaevC7eBkD37LDWX64/lOD7YdKG1o3yUNbO4tvQ
CBUIhzHKiqMjBHvj0n7zaXqWpaMhj2oLDte1lWBFXlCFj+M0r0Dxa72RBVaOMfbLdc5jwLFnIEzR
jgf0MwUA8chLwKcr8Z1L/g6jxmg4yv7MiabbmTyPE5YmHpuvcxUw3n6pEWwV//U9JJf3BLds3dQo
mI9g6hHKt00OrMSLceODL7WYgyAF/AveWyJ9dsZTOL2ePtDPkKxWZddbuqMPQHWxpWpwiQXni2nu
xmQdASjQ6kjTC4JueYLWMnY8IFTMpI2R0ZsArQ/HYaCCJdnxiZz/UTNXfghWdlNSJWMTotAMokn+
oG3WKQlAeQIQYlc8U6ulmkvx8PsqNZ/bl4Nti5yJ3o6Gd6QLmOiMGrSb3TbREjMwm2Eb0F1HO+Do
R5FwOhNNj0wpZbX7guo90/DMpMvEePuxKAVX9B8m+Kduk3FDZ1oIRKbeo4xLE/UdlU+Bi4RQS7Cy
qqUgTQ5egPkZENVhocYjVlhmfqJ3IWUnJ/aMnOgFqKRa7j9sf+9k1g1orZsB+dXn+UQtiHMjE625
4/LURj1luNpJN7NPayjE75011LUrdOzHwpYKspe7OYp0ABIcVojZcd/zCzRbRwROZLGt2TdabxOG
6/OtmAz/O0eYnka99XSoPKFzgF+wMdhnv9Jfm4X7UZMkhf+WqmnDnZVBjfBzPf7jPHgjojKVACO8
xgLZxgAoc96SeJebuVgO7nbHLM3H3fTU1kaXIhvDryEJNXe42QiU3B1B2KEKT4bGBtMIWI66Iwy0
rTAiMe+jo491zPdCnZCMC3iWLkBaLW45seWxRib/Ev7PICL1mJUhSZdEF8z9HyDxjbIQhXHQIKhV
UHvMcvcBs812isVnXbey5e88aUtZBtW/6KBhQAtl2/gJYkGbf1vTr75QAywpBkvTD0PSq5KxDnD+
QY5MOACi3xufFMNeoBTGlYke1AHyVmOMKrx2aIzxq58xYSkcmGDT0YPawms1yfcb5Gmok6Ul76mn
G7FjY10igRJFqTq1Js/9X+Z5cQoPFaeLj7kQSVzmwqEneI9j5kI13NMypIvOFY5mRevsH3ImW3e9
1DErrDIHOnHSiDx3y4ygO7JE2E0Z0YA1r91qzv0uxyynDDKMX++qjjaYhNt9kZyV5tUd+G+UC6cO
bnXcZtyzBJnmAqhTeWyA9PoGGM/mdJblwAK0gnMQStggYjG1gcgG15IZSEWTxTZxvM8yDI9iCbDn
QhO5xIS2m80tv4koueJ7npIlg5CjyPF7wskcZaDI0OXW50zLOuW1JE8re0IH39J+TjmEhlVkJUmI
M+MOkiqDCP4YlHQDrTAwiY+JlrdL3CZuarfP2MKKCkWVXq62vUNoqmy84ltkkRPrsrgvMthHKl6p
B5YR7EIKyWkvE4rxiF/0I4k+4RecC7wL+r4AFDLwOd8l3qPunx+q5ryNDWR17IZ8rO2v4IJxJuCX
BOck6GPni+oOHh5+K2vnE8vv8AuI4d6+1AiM+ZaofFtkAbIkTv5OGw4fleBg95C1WGu/qH9x3K52
zlYW69h0bAju0b+ENVEq3Thg2GqzvOS90YY15Iq0hxL2og/YgdoUEhC9/RWHdm4Bq5wJNqykkadK
7CGQqnP8qe7edjIKvc8Ri/3aaQLD6hN0l9XabeTOfLnBuTnPeAVOCjj5KINOaWvSGO2CyPK8i39p
zGHAaH8PMhsZniXsoSMnT4U1rMMiRsuR7ykOZpop86dxUUnsIX8aMBj11+eqMvSHtUwdQUiLJ/ua
iHYsuWnHzhuK1PRWGUNn7XBll0yCa2kBUMSpVrSvAyrTBlSVN7/OgF4Uh6lik5f+OdbXNZbNzYgb
j1gNDPjo9doxYSdp6GfOShfZEIDkbEsIlewTxu8vyiaJiwHM/+Pz2A4Dsm6ftYq83D29mgUh+2kJ
vzXj0LW86FQzdpVM2kxaDsEWPDCs5TvPXbfNbyFFFDufDVWQx4juTmGTCr++b3r4Pw9CTWyHap0D
a4KHrIsPpe/clQzss9To7/DoKiqTkG3cFWwSkDCaOSvOo8J1FHRZScLrhcfb3WDZU78Xm/rSqZ9L
tcH6itQ0hgiCWrT0tuvpqm7Wd7/+oginNxnWmRTxkZXKB3wlLauA4skYfYWFyyGPgjzgA3RpKqv3
1Cn9fiiMRtwCzcS+pyaiiykYI1pKBQU64+1NzgnGZAr9ZbBYsixdJ3tJtke0g5F9TnDS/JL6hRl0
h17HO1AuiUaMAap+wfyupgfHro6kT5o2l2RTp746542mmmsDQWf108EmljViDPPrDZrF66Rt4mEd
VKynSG5ttc8plagAmUxIkTjxOsB59YEF1j1LsQ+h5EhUvU0UT/lQ0o8Kbr2ZWL++4RtYeJKSPOUL
Z3I50g4HehN55y+ZRCrFzMXnbby879IyiHVMmxfAsgwqEZA1kSPIqVvn5BHTv1r8tT6syciv9KAX
rK/MOpWvcOwQC9HOZSiMc/pS0kw+ggG77LDiwLnvb3v3SXDvr3oemLjoKAbNv29ocIT8g39xhpp3
TFtSXCPH9R/T378C/9jkHSm1MCOXdHS4gdUh5940kMTotGSnUOXp0QRwXLQewKzBinzskJ0ITFgD
NiD49PYA/5Ps8nOg+azF2zLeKeHOp/07JJRKSr694Q3gHgDlGLg+A+oRUr6UaFTrnxfmhDRiEyzy
afWoJ2864pGcF8JVAoin3vGALTjcXG6CeGrPjRsxcNf6Er3UDakRklSSEbEBgvCaikMi03nJJXNd
QkItRutJn0cWchiuCtnOseLOEBmhZQiCoCUl77VnuYlkFMQofzlxbkME02plwgKcPGFonSF5Jmvx
BYA9o7OU0EXg3l6LmGMZ7UfIgn/huGk/jHZDWNBU5tyLwE10Pwu7QUSX7t1SXGOMcpIK5yfSfe5j
c5QC9rOQvDzbJ0xzFATgOqzdKW+kryN6I5Op04wIdx6i3RvaoH1LilC+Suqxq6HQPgxKElZmJTt0
hfd/O5/Y8SWdkuhFmKI4xEkkxLrnwzd7+MzK1oBnxp4jULjRBUGGAw5GXp3wwhgAtcUskMXclaKB
Rh9UyzCC7/+Fy73KRXRl7aPHSMgvRp+CvOvXlpnPwZuYbelB/GxJKK9Zw+LM2gztrk342hGe6+po
wQuyGKVGo1JHcu0Q7FuHDZTRSUYST1FpeapPp/m0lysCZ8cStMRw7kPFx4LtLlp/zdCNCJb0HatI
LgGR/A8YaIZFtObGVTfAxwGuV56ep9fsvSKSgp5wK60ihHEHSNpOcPy8F/T/eFx1GVPeFvdmfQto
zvSdhhE7UN7OrQriITXy0Tjq3wsoRD+EjeIId+xmjpW9K/0eCAKMJIESiVaWgcf6y2I5mRE3oeTT
WI/ouNJ5mt4uZX1aTGur2ZkdS5cUpcEcokqbHW7w38uE/7Hp79RL0LK/8SyaE6cJQu4Nwt29lJmj
CpNhqPhDdSQDl3RI/ykhB04s5Z4gPVdi8qpQwlaxLzZEk6dHXpD4XhceFFDdLp56xzWjXnV7zBWs
lYcg29Cn1YCGMFIiXfWumEWJ72KP5uvXFoCLpK1gbYAb78Zm6A1D7o60gtAXasBb0TdQ4YZiQZQG
uWOpDqJsexLA11R9QBLctLwBOX2E00tFTRnnY4AfaKq3oamFZwweS1a4ZP/cEL0idOHzVOPJ2WH6
ZFtRy9BpR7qxTqnn7ejx1gqrIeo8huqqBOWgS9ZettlnnBKCOq7mKUC1Ly7lj2AhTcrGpEXJbNEo
7c3g2M7CkHXDcZ2Ol0z7v+fmu0ieTz1CjdJ/9TMuWVB+tR7bdbk994Bghrnx+EWSvUM9csY0460f
9nEbjLf/v+AVjkmLULEa7VRjJHjV/+W1EQ0g3mo1L4rG+QejukYd27iDYRuEkBLrPI10RzfK6a+3
OutnGM6ei4QWeyaLjf4MIZnZu/SujNzoRbLlU0vCliAOOi/5OPKO8ei/8xzdt99PNPiFB52WxQgt
BSEXkN+yBx2Lv+og3LrxB8giGXBfU3R4Dl3+Q6QDGqT8gwf46EVIwEaJ7aa5qOQgQZej2ar5aOwO
6zr5a4lgPrConfSggk1friirqkmykRye9/UTY8a7zLPThQVm2PI8yL20pYNkzYrJtbOsI717Te7s
hm5T32sF1d2XM/RBKM/ESBtonJW6tby+WyaEN407haSNFQRyw9pByKWadWpCxvXT2LRMwTH6RD4M
A2a6HuKaSWDquHfGWmE4nOMuprzHUWSXOBribFpzh5k2nsedMtGT1aCBLnC02Za18KhFBfdPyZJP
X5antZy2pbE6kZ6pDIyoEozDELAsPwcdpL8GVJAEXAec4ByrQGunaaPqUQ5m6zpo/CPxwPtHe6/P
KRiwRhCwvOnAQGbB6Jdl0/L6NWCYlyG7mVR1LitZ4zc+tUMlfFRo0XnliQ6AxBwPP0JnTS/ectbg
vW2j/Iekjg68gZh2dHcMt/KEYalw57i3kbuDDIn8bMXTAL8yf64eK3d8b887UxkBhO7ww5sVoIyM
rPHGHLntsgDqdPuCeg1JjdZDrlEXIPmhGpl6aV25y8Mn7NzZF1Ck/61YomvX895di+0w43mZLp9F
H8onysb1Bq92e/cD9QccDdg8XYoI0FYV0ssOEysO1ERDK+sXhSX2RBlzGE8mCbPFYiQFrZnhh0VY
OL4sjSYA6vrjC5PHhMBiyKwQ9muZIL0zhrFSRDH451o89nYKmUXro/6EaRzzwlt96cjML6DYCe7U
JMBYBy4p61FWACsOYImfzQvYYLAX4O9EGyf/ULDBBlXZ7V44bR8TjPTdS76105OQY+/sjoERfj8C
ZCMaj4eL7gyShBdsU9b7DVjva1h6V6U3A3yN2LW6B9S9p9Q7+FoJ37e6vcQ7ZS926mMz3RJm1bqj
M3PbqqpbgNS7j7R4XvelAj7Ci3GEybyEkljQ2yFmYNrHtdglASQqCO+yDmK0VC1nlVXcH86UwoOB
DemVTfLZB4vt7klMh2oXfATq+K1unhEHBm33vHqfubMsvvz3CyOsDrEg3Ya9K9OZ5IRweDD8bC1g
pyz5kOJE9BiKPYxoPDmMTwtY/tqQl09JDdzcFg7kFvKyJao1kTjw4QOMgjiaWSkw8YKL9Q+CtWC2
DebAmTgSAhz8YW+1QPvAr9GWxZfWnqWY7v9V4O43OZfpYKqQXKqou9erjwdqQLHSkfdEH/B4a/lT
v2KzEh8xLMJ2vj9ThzGm2gEXtUOokC6uXbwqS4QDkpCcHukSSFYjOmOL97wSJz3eHyrp9fxBe++5
8An9+wvE9pWaJ/+eoInrvvy2dX1tghSyVhG2Xga9pXoiTTqvDB7q82dZBh4m9gsew8mP3I2snj2S
7bGk3FIClxpEyJ8M5ERR0e6eJ3MvDWpERROF7FXEaC4mz4CgB5+PaHlHbcYoMhGK1gO88lY5CDV4
huaDgfl8MW6/Fbt2oZNApDGcBIE9XD9RZoO97cmwtikGRatBbM7/pnOBdd+QrTgtgxEQweVW1aeF
gNuHQva+dN/ldNzNXf2z25pKlpuEbNomojc6qH1v0rn9WkVtFpH9XX7MlgYt8pMhh/seypb+TCzj
R7TKsd+nSalHOovyDXeWBAqexBKNVpDTNUGp0M97EIkDWvCXQBsUqdr3i5r2ktkWc/wUmhyYwBNF
0SQMPP/CanmbLEPeOMYmy0Yx2MAD5iwC549bCotg6J+ENvDTBuje6AMaiDWK5Z5NOrOutH2TGiyG
xSX+XX2I/1uINILn2c78Wvyt8EuQRRx4d98Zeouqm6YxTWOHe+S37sohTwtiYosdMa99fmU1KirO
TC9oHbyz8gzwSoScbJOzwgjBr3iNSNAildNVlmoDezkvZ0wyAhLf9pgkrxMSYnYedZxnenfp8FA5
eldQVVTLAik08YY9XSc4CMlR7ldsAU1ZwrmNf7jILqXvp4TWG0lw/30RpzUaMtl4Xmh4qIOUMdk9
mub10nSLydAiRmIE7oH6e/Eyq+jcvbgxpyJI4McWsCWxbxGJ/3jX/rsTucItNAIz4ZP0bsZJ5zUs
kULFWLczzkxGuYGGGgZ6E4CYSau8oJpm5x/hcNIV33xgQdSuFMfdZzkwVN0/c5jDcJAh7MJLVAUg
HW0tBPT6AZ4qqfMDf7chovyfWTMnXaj6TmwjJQG0sKpzZrQv3ZnJfwrwMPEVVwukzuyHo/z+aPwe
MGV0RjEEy03UeO7VJ4I5hqQwfdqs66URuqMZmnQqWedxXgYLOPiwjWAYuShQyDI8H7U9QlmJx55U
EuacMwCe1O4IEfcqUpbB4Ua6KUVKMjRFmdQputQ7rYKEopKQsD67N0+KS0MC/dx7VnVj1htRUxWN
Ho4HxqCC+B8x5Xx7JGHk7X3Q4fT5OrkSr273xCTz7PSEbw/mS4MhmghNB3OoQq1xztAf3htdg8oh
KZZNhS7IXuYC87X49Rg1rKciNaf964RdbZyR66e+AWF/NYlzmjkdwJvIRAiBSKZwuwraTTe+WBn1
DekQCnTBS4nQ6GPhIeD+cNQOgovlevpOLfWTf9J7LCMeSTQY8bN4gPs1Me8pQZqqI540mQFrbjA9
WT9TyulmspjOR+qnm1Bx4JLUydyC4entMZL3IDt75AK4sBe6IGTSNLzavyTWhJ//VozkxBfuIbkF
MjlBr3Rczfp5l//sI/tJx5KFF/hpp2fr0bOvGyLDNfvf+7cwGp+pemP1YnaELnES6PejHINLSRI6
lQFA84r6Q171EHKqNzcsMNPpq5X2Xi5m8ubNzXWS69n2CzO4Rl7GJtziKdIg/zXXVcy73SxyoLOk
O4MIwNi3lDMAy9Xbba2H3T77U+Umm93IzGZIhXIC/hG1mGZcf8xpr+lCyDgJvpJaEMDJBm9KMyc8
pPv/oOlFob/t+cZJlC/naq8tLCLzAZHu3xjR9xj4aWLm6j72ihI88NnkHYJ2gGHPr/D5Y+3aHNs3
04EUo1p88L0YRrwrpAbI/9Kzof4uYnVS5Z4Psxeep696drsx6Z2SuCpkmsm67vehz9tDSYCmAcHq
ncfiCX5Sjb0V2hBzwqx0Tyx5OrUDoKpZuJUoZXc3IKYVVtNg4l17CcsJxNrDe/uXVwY7X1ESAjDg
/coNze8HyHjleEV4Cx/LNXgnAV/bu7vn8yjqycSeqLe3IWSHD3JWa/LlCAhaeZt7w2z5h0COZdpw
cYeT3YK6ivZoJGLe7vc0PVMN246zab17oxD7nYxeS9Vvw/HTwuEGIfOFqJa8UJoefBal/l5F9cOI
UccmXnqtSobgEBgRhqWD7UlZMshTJ8ypTj37lHqrgVXJOsaMAnRKQuBVrPCTMFWOAxfJKUX2nr2A
o8Eh+sZc4PO89PcYfEXvcmHhNvtzsWH3MHlu4lBW6qbXy3gUXWHGBXaJ8X2rgZrD5rVChL7d2uzK
EjN2nt62HTsgkQ3JUv8ENql5PVGt3+fFO8lO0XACQbTHEIhZWjYcVWMetRV8geFq4QzyoprYaXNq
M/de9uEzKWML/P8IBkOiwopUmBuaNQEFj5STrqpql2m6jk+0ISwLmDPaNfpY2eNlC3CJQMnUlR91
fnCrBw/WoEllaQJ0lS2QannZoi/AdwSrlCm1V25k9/N/cyObsJjADUefnO2wYklj4XOC2DZuBDZF
EOjjzJqxjGYSRU0xReC/mio1nCCX9B6lUuJtQD728OGxqFNnlXds0Y5mmMTt15DfjjJBeP6qTx4j
eAABo1g07yfm8rT6nYqFoVIzNlA/hBDmvCLOmljnOBpx3LQSz2NhX0rwfjCTvl0Z4yNDOIDYzyH8
w6oLsmR0m0DA2kwOsJ1w5kjC36NNiGG1S4FpV4KQM3AGO8RPz/glXde0RN8kC68UTXF2UhWX3Uog
f8dxiLQcQFc3xc0bZhI2YmWvN4jssbwLOjKYSnBEZWdZFYdM0c79mWOrD1E6gXvJosjZKANhzPfM
dKsWgV4bFy+ptbLjI0anddzhF7e0YSkEcCxowtjIrrE58Ktq/6qgJMHyCz3jMNYD0lYy0Gw3S0pg
yTvxw4il77n17utIV3eBHsIqTitHaf1sUn4DNcvuBcYXZgrccun1y3hXv/b9zamfIbS3vSCofaKo
e3qU2gPHvgb/cNAboWYh2ZDzEMbCYgehIG6kVBYAh6RNTMgAw6rqpkXAziKWy2IzvxsmHGBz2RjJ
vK9bPrKS8DkSHN2d/GvwhXuUmd3YFBV9IK+fsFtiJ6KIpCFngCW2guCJHhSahR0ps7nme58fRcZu
KHVi69JTncfmaRl7mgrEfr6ez0YNUmHw4L1HyZ5tR1M6CGaigh/oKX+ugotWZ4FbhQ7nLgWmFG+3
dAue8wwvxojqlseM3AGMBl3kyTuoQTaUI1I4oUs1k0nvQm84V2nx98MMTFM5Uzt28mNLJ7WfnfUI
Msd78HzXzoFVu+7fxe7Hx9wIygvu+qeM71LP0xNoSfp9JbYzQpjeoQ81qIAvEtXYcuyZSXih2pV+
mfVPtjGpMu4T685UwcdBjLcY0wVcHb0A7DcXQhbjNU8fh9ZEBii61j2fJRTTdHuEpo47UmhdSUgS
1lcRCqOb1qT+kQUMSAk1DKTk95TnLCpSBfY+W8GTgFBIhXcsSzBvbQZQUEisjnqr4kWz1vXgnCqt
o/AZRIurwOnp0X6nWPkJiGqphZFUJUw77G0fESLoCQuTao2qdqIhoIDTOCAxIXv6phhUimgmPS9F
sWY7kk5+HRZi6auPgmplxERAq1XAXKgmwCKF8PYXtxaHnGdo1T6PQ95C3nnu7IemiBrJMFiPvocA
ly4qcqmXA3H5fm0HU55FsnwsShwlhD6WIvWYZxtYjTdI+S0l9qAdzOyIXEo9amfqQDT9i6KnUpm3
wGEe0YHqVSE2do+9Xl3dh9ciPXSV3oOl0mjWaTmDg/xsd280rwF6jiqUaS4EJ1SKz1Cy5Qbj7lKE
XbCxq0IsRl+7Sba7FIUez65vdd84ljd+y7lfIUZ33Sr/xj5vPYFc8yFIHeqOJIvchANv+3VcQ6To
FU0kGvFXiej4bLVzAGOVUthSMKKQcY7ZRcnuDxePLS6HjH4wYJbbJDqH/r9y2hxU/A86zaaHs+uV
q8c+sjULSbK8z3UCX0KYaVxGuozSGTflWinbGeRpftcriX6KKhGRZP53RZT8QQMmeZRhee0SfTEy
NErGyFA9xbOzsOAHStQY+O8Anu0lP37FdN4YSajQjSgLuj2t6EhwKVAnBjZoDwrcqsOkBucVT2Vu
/mnuvWa9GG17JLAiar4Y27tmvrQThjB4PHckHL2DWTvTwMpcm3TvjkTuHa4HD1qZfeNUxSa7cg8n
qX31UM7CPwK/ZxuswXW80q/aHApDFVLyYX3FWk1/6cSAdcFxUJdhkyTDzO8kN9Q+cuGCpm6UKxT/
aay05f7zvcgjlgAOxLbjsBdDtST5gS0PeFmcFiO1lSp5x5bbBnFgwOt/gIjEYXgoYqdeqAqRYMuK
GmJNlrvFjfW7bQRqe8QD7qRl0dgVhMMp6jDU/Xc+k+XyJcbbr2SAWzautuuY5eI8EvYfO0toH6Sf
ereIrlwAhy91sdwfaAtEojm7zgSvY72Cp7iqykXpV7jitoIt4eLGEaFOVCT/7zIfeqvaAwbBTTkk
91EEOcUXQLxP2fP6UlCFPNL/a5viIfuvglR6RGNM/b4QB6padNyoRnxRfz7LDGYpK8/oyL3paUNV
F4RXHSS3xI2vI6ESomsJjJM1SjDADm4XJrDCcI0MV8vH2tjTMTqxbGVuwGU0pcVSp6Npq4sQh8tr
O79gh3iGzaPy00aDTxv7yWODo6qTtupWXR8FVDMtaPM2HYAVRDPI9VGXjYsd/nAoLH3mbNsnPvmv
uxMLODSRj2/JVMmE2+kyZIqiqlXZQkG2dRxLsalYKd1xfuDuNzhgPIA0Nd9hKk+N2yh+U+kQytVB
mTxn2NM1ldbUqgflQ+qyh7JpFXjAYi7n53SGPqz3DVgdNLVDz5hLARd8X2/UfvAoseY7VJmHK4/B
p65Lzm64bcl9RPcIDBuJvJpWsI7BibcNFzd4Xvzwa9qIrKIQzmbpIxdFLRoIPlFf+T9njwpIO++/
SKBQ6kJCkt8kUVIU6PSRfNHRPRxTZflswfomIm5bmzHhnS4OWmFQk+Uw4QdQ4SMSaRjtRX3KQxdS
W0ES1/MAYlVc/APw5FbQAcLOLPhzFhR6lTk3lkbofYJeC4gCZZ7baXbgOew31+dfFVHg/ttuqGea
Z9IDb7fRUBT6VisqgkQ2eAm+XwvlJ74tFnxsyvwlQ4W4tNsJXAu0aBsrLYg6IJ0P+H3LUa3Ghxj9
YrXTE+DzThe1/Kgul2yX6OsDaSAe288LTq6uiq1NvYm4N+vLvM4W518EhpUr2UVqZG1/Nl4fqIy1
zWh34lcaXYnO1+BOhwxIvT1dvCGmS9GC+hmviGQQhf+gfXVbosURha3jnGU7rbmqyUbxTpP8Ch4R
ZV10jFrb0AZSMEcOyfzKSkWCBgGcf+uI3SJ76cwQ0sMkuVLxFSDp0jwmdmefrmdDKIdWowui+dc5
0Nd6IbeRtHRj0VDWNHPfJzU5JgZIV0JjE95/qi7H7qtjuUKy2lbf7WtsBd1poPEn8da+kz9yRC51
E7kK1spsEiMSzFucqcaP7LDtqltw7vuxJJGBChVIIgc7RvdfsSm9Ss+aT6TtfpmvlnWJBqD5eDb9
/IR8GBtVcOrZZlaz+g3GUXLdPR5rV+x2dXw51NnN1l9251igzWPv6ix3jHWPt5PMbR+DqX6u/dgi
dm16tFgIBWy7CY/Iy8d1JGm7XDPakfazSitVb0yWANH/h8/swrGkG2wAeuesL8EP/+ZlOYQ6xOUt
pi1FZdtaDJrxIAwRMRl4eGuMHsvpN3WpoYDDHjK7Z8FIJ5Zq2IKbfxUkYRUnZeRxcytEhtIeeCJa
Td+DDXf8APxXPz0sHI8K0VPiL0eZm7mBFeE1pnhrroJReG2qkBhxZDxcAFp328y8n9miO1CtVf3j
QyVAtIPsheH3THBWX0BUaHRRRrhdSg82JbmC3OsQzuEjdaKNy1EoEJcuKDPhmVtZbSsqH6gIveaP
iqnKyaQ/2cOreC+gsxSsCZ+ronTLEM2g+wB0F5zy1uUhpvDo4O1v9K3v6/cJRy2cGRVQMkOoXTVA
s6ZKMJlnlrI1hM9H2F0Q6jn3hVGldz2ufLnOfYxrSgo/FkwXKRtGYOmVJWFsDfKS12n9lHyQbfSW
PMxr5762Cty03GhgdBAqWc3EEAH7/pVtIIwsdxeIZSYFxpFaXhBg5tvfBHXojNQ+iYHHB7bvhrYa
+Y+0+mYHPgMeAR3C7G8R5GD/i81sDcU79SFFKRNn3jn8Tf1FD872D1BLH5LS1DRnHTVzMSmGDlf3
DYsDWLlfjH4l47LH6G+aVmvXTSokJ9mOZHl8+1BGmnoYAw8ulWkLtMCW4zilx/C0NTRXlA9ci1iz
CTArEetnaQuvlembxVD1RxU2a20/W70kJGjdvmJX8DKJbZyKdlEq9INf1pTWrGbf0IZzmmQMbLGn
0Ynvb2635zDeNhAZ2fiCL+He+RFCtcvJ6+z/TouqR+dVoa2N6q4kzrSEeUO6oGWznwWsOwNLsBZx
7KLMGV7Da5u5aECDdL7Mao3c20MCdk+GDsEsb6JDPkkoY3TPGIXcC9ALNn43wfrijjcuB4cJ0/Fz
tyoAijE2+gNFR0bQWNaFmkkyK3L681DdOYMHhMGLbVU85sP98JXqQfjoV/KEJPxD7ltWoQvETWkU
OLRQLlt0+JQLo7LACkdDPtXk4AmrFZUSh4TS69PlwJ2Ci71KCp2eFCfINqf4s3UbK2nJers9DzGP
cyt7b2TWs6wg6Y6tJlNDd1CSUlsDj3Qv6XJuGFJ4UjpYW30JyzxO5AE5IyRpmxNrTYjs3q8M3KGC
X0dgI5ZtaH5RbkoquANBtO+aDcGsJT4guUH45uOX5P9174yjO8380+LJ63bY8cVXbrE/3+2QBATv
REjQ6lXdvClFbIhQ7/naL7XZXNk1rxBa+pc5VwbNZRUPtkPTKE/8aqcfUZ1JZ1iJZx/nxSuHnamL
0PW6Po1oiqPslSPURG91FZWmB1EAmeRGpFeNjoW5TM4RWfIBe6IyWbhFypQN7TyIt2NrAdlFxsVq
mN66ZqW+NV3C73wQSXBOwFw+FseiDvKGKiTYa42cbdXqhcEl7hRueDM7txDkhEbJKk6lZI/FdkvQ
WREH6lr6zDbeK2gyACFjW6aup3XkjHhWUGTsHQR5DI/2NaFpWtVsc09k8V318wLUBBoMGGzcwF2E
rApJKxLoAiLP1xqeSggKVo2cgmx0ZftvQzgQxiqQn1g4KzUkznGPsNh4OXd2yI3cb8b9Vtivpvgi
oHab6HE9NHlZXVd4jqFwme+5h3Hv3oNa5xF5aEGfu6MOGspaxV2z+dvcJnrvBtCKcqwU91TpZPFU
nuSKoi5Io3fJvw7jtbbZlHz6Da9nPoGpR5CMJGeQ02C1vvQotIcwKUrU37dHs3rO1i053cCUoFGU
uBNVnKibXoz4zqzFRuWUNKOxUXVoPafYXzr0ZB1XFm50TTGACflKKrxL8imKqCgaFkL+lO5e3b4h
8ayc0ez8QU5YIvgZXQpgh2TokCV2RSgQsZE7Td0ED/Zf3DCW0VJQm8H6IJMBiyEhAJukZ6Mb4U3O
N880SM7vxNF2WyAsShrNE4ai1xwKETB4IleFdIKOgLjmEC8tZim9rUcIe4VFLFJszvf0DFUzoBZm
ko2csZWT3KDOexYtydan97I20KmDDYGyPneKBJqWFK/IZ9KpQ+B3GJWQF1p73ijAmhQxQuBcT+F4
rjfXMHOdaAm2h3qGc40vKRZ7xEL0dmv76mau3IPAGd29sfvDuK8kLhyplfA/rVfhqODI1s78jdhE
yi7/V4CssBehjIqmTrDSNsWkbyUWJFkaH+vwLWI1YEWOvwtiYnlzJf6TwFuax+/ZbfOPJI60pcMT
Sng6vcU0MhVvC2QwX4hLmS5g7SoiTNJe7m1DP3u/FhDgWFfzrmJ5iN7/fQ5UmMqGeiHOIlWWDaul
tra97zA01Fwz/LbrcLTjLZ10C56sq4KIluJjNA79gpUqdUxb9uxOHDdFZurWL8AUovHg0YCsd0wa
GcKZQi/+7/juDIXkTeW5wELlumIx1VGy6+NkVqKHAG3fHzAuFth2JZBz3xnTtirwkhEEZemRVyUe
5zevTgjft2quZ6/g6ZHqOE1Tc/kmYsq5THj5t5xuBshe53vQ6yc772ldwN7l74aV+beZLd+PjIFO
1G1+fqG+uGPLFd/abcUxHsvzcY0LatecOMdL4IzgExjDvGIU8uy/+7CQ2UPF8Knc8ksqaPhumpZo
O26CKIeh/jJ/OACmZnrg6q6CkKJCgPgim8RepxjrRao41b9UfJDXZRD8Tx2qiwkACiKLV0bHy+Hq
9B2jF19ErFeDVn5zMsJyJ+SxSVT+P2SHi+/60Pbq/0OzP6zrYxwxhz9jdUOwDKXugik3NHkzCuro
++sjRctjT43UnHQnauZnXx+CXLF53ATQYNaOzVgHFhBR6pDOnjeRR92A1KYM0X/6l8j7ceD9RNtD
S+1aimPMs2792tv5oVmWOplVv1HPIQe6UV/avzJlAHA9B77nLL7eHuu1WiOzufFuFASFF+2FUn2I
vkpjjuhDkRgZAoBKc1/bOh/WypUanq5hyecnI1JbPUspkF5MB+qVFrqmUZ4dakGxM0yvUg2b3pMV
g7bSx+xjrZCTKjEscwzcfzIkhjoGTvL4V3iKC2IFBcnsZDTBP/iXZSaCT1ryaNJM+Ub8Ij0cl3p0
VE7mKhQecrQcTKIziR6KzUeYnicnMUSMNyTTWty6xI8wtIcJ402rkfs7OfhhhqFK5IEo3NavUhH+
Iuu8+BY0cEF8P3HvX6I8GuX6xvFStWnnB6/Racjut8J7GlfvXhal93B6j8SwwWTReBQ8zvYdwNVe
mNirDUC9qGJn2QC+lOdkinqd+spifVm7qBPujaU5jOB42l4MG7JVX5M0iPSq9jSHSD80KPuK3+ek
83+ic+NUdSHDsPkfca7W1L56HjXoeiVPbvm7I0qNd3aYvtttHFPijh+YGhb0lTnm3SSv/CBzaWpI
63d1YLLKI+AXJdVyr0ceVQxrnY4F5Om03KGZ13PI5Hg5Lu5n6+MKE0bSlP20vGiFMJJyTo+bbCvF
1zXLOKIl+8hS96esdlTUGG2ZNGA6gaxFC55QyiFYqQwJLDg1hNpoDzhMYm9r0jLwybcel8abm5BF
IYe8r/SeLz2DaiekptFos3VZWa14mhKCM8p7UdgZOcYbVqeKLKck8sScgXXNHN5ilvjz+KBrFD1Q
jG8E7WY0p58XQw3KC8wMRrLo+AGIVdkzerjX23/y0E0G5H8/juZFlNNLeO+4pI43aga7fGrFak1w
FPxjDhv2jckLD5KAyMRSPcAkYlWQ+SwMEkhcb74O25TCieP2TevSxs8uFeqcuWikjVYPl/YYZngx
/ir5bqPtB7ADpac2XvusaJhqUQluUINInL1LNYMC858bk/0M3HlHFENFCbkaXgHkYDSDSWjd4O8C
ifZge7EWWcEExb8JtuB+ibE6c4JOvwOX6m+PKAIuBhxlsSkLdL+4JyxmEMC5e+ZPDU+L/PcRPTdl
RArHhlh0GV9AXYTf4rxyba+j3TwiHSOZPAmTVGqNgSIYKdjfpFXzJXjNPXv4OUl99VLnO9NsCVnJ
f5g6/NiMjlEBE28D66SSvP/jEZrXA2hRXrJn7RT95qc4MS2RLK4vIK3nQaq0RDQmUCea4TqEzTPy
L7WUh7wlSaa3sNTg0H3jD8gC20Ko1sG6wJcVDRFbElBAisUb3MjqrgGuKK2kJq5w8Ne1ZfYkVPYo
jaX7Arkk+MkU46BriU4Jwd8jF6O3kayaJw6kYJzdtbf1mDGBq27dyWlqsa/Dd9xGDFv5Z+9ZNddl
37kZwjNgRt5bXbXcPWNzxYVN+a+WBej9fa1TEP1wOCBx9AoLrQ/cGWPLXMbJK3YnYiBjfsu8ziuv
WohE6Icr4MOYZy6BIKufRaiHsxRK8waVmBt9jK9qvuGEISh2WMitNpMNQNpaWDrkja9M9bksfnTd
ydBk3PLJMSrUq4n4iOtWu9Ev3c7woOD0ree+eNGXJb5wJh70wNh2iwUlumz77C/pbkDXbOT+xqkg
59pAe6pAFSjnVAaG23e0HfkWagt/0S7gqdgBlQWA0anf3htVYU0g/th+JhjkYpfdEZmaa7fLbjID
5S65QqBapU6FjWDCBt0WB8ZPNaaC/gRzgIvitLEuWyGti08/zYdRADmsCu3Spp7cL5l4Rw3FdCb7
CSYkld30kD7KZGdXmX3/7T7je/Bf6VzdxblCf0otXYUj/1y3oAurS5NNdX7AzDRuHLSAQ3BqR/Ek
7q1e8tKMTm8p24eoz29wRIcp4C3ivrFyhOgXZdb68Ek8bBpCmiwkWdvLUIi9MOxd/y+JKqNWn1oh
0FydenQt3bcIPGfXUw7kXDR3k0oCgvqfzPTnTjOkz10uEZuUKBvnabVnI9OYJwLKHsBzQiQd6rJM
2wYSqKkmUbcmnuAsaeiYUwS7GA9UcwTscVVY4uf6G85EEsGF1WPG5rp1FI9cRLlMH5yziCZfY0o1
qJQzOoSkziunWKifnDyDoxLwdSLXbF0HUKvZl9RQ4ZaLzVvZ1lZDU74RZDAgqNajkPnrEmnpDK28
4i47Ro7NRBMed3/Qn6y/UMCZm3KoZ33V8AthHXy30bLSpwAAKSMvRGCHGZjcjBsFbaOA8/cMdv7+
OEOSftUVh992PkC/VisW7LeM+QY4fg5xZTuJ3Q+EXaCqWIU9HMd8dW7aUUphPO7uzgDYoeoBvLjX
+bhCyYNzN0h+5dbu3adu1VLqDTu+xwNSrEHyr8Cc6cGbusqds8nC+QrkTWOAim2+kYilSZrbn5nm
EAea9wptsHqFuz+EDu0oILFFzx7G6GZE3xgLo9EQ0adbAJ8ooNYNNHjId4iw4oi+b6stjUvphZO8
UPPwao71+nmRsxJcnMYXyVV/IdT7SucbiAl9tBEhYSVR6AzO3NZ49RM9bSOg+TD0g9mtZuK5BC9g
EwF9hIw8vQiB9nlTjc/LygvFoiea5RETaqe5QtY/crhd9sJmzMJonJ040ochE1HE6B8QgLz/h+uV
fEeDjql8g1XVyWzcBNSVYcxJoREAHkQtaR8WrQc8QUmIUb0PPad844APNx4Ft/+n471dXarJGC2W
t9MXZ8QFPh+egsI3vvlZP6cB/wGrCCX0ZnJBjRcInszwWlHblxH1u/DR44GS5+jY36c+JmGS4kl7
a4D2NP1C370q2jqoAYatepcTMr70oo/9u2kAIHEIzErJzfBIX46syt/h51JN/QfxbcZwgfZBrtbF
zLHtw6gKoz92tAwObd3VJmBkF2CoXBbi12kbnwyqi+FNIRC3O3MSOiB/Z7QtmsXcPDSJHERQ2tQH
uE2EPHrTsQ4W5Xjvc9uBwXQG3P7yKUmu5ZXJt4cjWeg2h1QFNwki+eVzUqMdcgAkysokeWsWlOpx
6u1IsNKClYXhF422hMyiGOTi5tQwRWx6ovr+hxt//1ffVavWX0tWulHSZXYuHJxJ3EVr8qEglJTX
CnV/de9mb9TwQlC3Ecs8T5QXDw82d2mqO3YfNNai0JjzEnPaFhic3qkaHlQGDKEQlPfJ8AcgBFyO
TJV0YuWOyJr3GeKxK6RGdZFXk/Huzm7RWeN0i4/6W25PMNn4y/YRFbyxbPL88CsFQnbWEsITCldz
GRXOkxjrfWxy1QnCjr8CwGPP2igpmADyNNchln8v/T5GjSdCsPrvb2fSWkiJnmvezO4aJS0AF6Pu
zeHG1lqc3F8tnbG9aGdnGlep1evlPr/vLV+TlTiDD4zjfNJZWzqpCTVmnmkjdXUmqd8r78VlQvba
8isEIexnulQdxlCUgPf7a6R2/eDqo2yG95+JfNOz2UtYJ7+0ic2W+XnzZDKZsriOcyZm6Q3D3TPB
cB9yC6i6DphNPPsup3zmL4/f8CErt1H63nUVaqVgFGJtccmFFrm/d+/zRCngaMupCkyQ34p5At8w
UFEqNF472ggoaS1yPqV4fKIagx+0wabTfOfPkPVMK4atuaIgvPjzAQeOLcqcmZluQt3ubBBwyMWC
APrcXSTFgjgVBQdHVe5qmFhPTTctcQG+AbeLonUs8jkI09jYXnv5YKB4KTX+NwQGOqJ2UgyYxZk9
k9mbnbEqBtB/5BTNwWmVMmP+oPxkuYsl1PYuTqI59+apSSKZitQ9P+bJSwouXxtq6SSbwgbSYZ9r
0r+yCBOyqRZscvIzemue84stH/8O19mJsWDY4t04814rE9UsC3Yb/2K3Pk/TapY5G08qimfIV5P+
6D99D7Et3GAzZkbOnCxknIzwY1RVe4otH7rX3QTQtISz83Z3v0zABn6QzWCkoRoDcgYibMMioyek
fBl9+VqVQHCeXbbSOdQyA5sxkuGNH2eik0gzNb1QdBEEd3Ca9iWWB1KuuDCwbRY5h+FbMPS65+6U
mWnOFJHS8eUpzz0TNi4572CRQ0IbLNh+Ujy3cCTcUSohX0zXwBFgmhjdxolvyCmzcz3HHhoxd/wK
87SfHArm99rhp88AFAu5AwgkOXB8jlwHvoE+OZpHeRdpMoIBAlcPk83f0Wd+9FnZGkFVa3k5uxvc
S9ZUQNk07RzoWtjX2/0kr885Orij8krRkzWqJVIaZh2jOyxUqSkG9TmD2vGVO4UwUi/0l9KPfa9G
RZcOUHpyUmxF4KXyezP86l/WuTzxTCYiUqTNm67gYAvrBpkMvCV+OkVONd37OnQgBOdk21oWQ+AA
5Y2HFv5nYAA1X/I2MT4E7zI0HLnFN9NlzKhIpgDAIds//kpwe1ZMAIcB3b1hFw03P2I5qDAlHRA9
UwWjeKKyx/JN0HVhI8oV0/lUgmWQLtQR91Bsw3ZvwAzIcj20wYH4N3HSsTf+KRXiFlAifu89d/nw
b7yHFfi/4sjjhA82PkX+tG+mNQVQgPuAayI6xe/cP/IA2rRSCatLYB9b2fk3geu5ufOHzKbzPF/V
Ls5yifuqKKSvVuE/tWou1uy/E6GEP4IEXO9LYTsb6zxAIXoLFiwKZJbFVzqv7f2a5VJTwY6w5Nu1
H0vIGJxiQxQTf3p00jRMwtdi5Qk/MErKfMj3Tz06PMEgmDV4rWbOI6S/QwCFK06GvLCuw7KCEx85
Egz/iz4uiJEiy6EVu1e/SL7eHTr7jUBgFNpHK8zB5bZGUSYj/r3KjpBLHqLjnvcNCD8Orse6QmET
vS6eGnaABWQcOmyVksALHeaqksq6rDAhRUwAfbzsaRlnhDh87p+HOHr4xsPdSmwOhHSN1btnN0U/
nJT6tpIuVLs4tVb7/hlM6qGlIamUYzOs8EfTKQGbduh6aHyZSKYOwFD6xntAt54TCPjHaKZAhwZZ
uyOA0qoxZCW9DG9GnWZsR+1lkbokI5YlNFwqRvfBfOG/UZd1xVLG3T6ywE/uZ2mwJIf6j7zoDeYX
MStc5Ixzk171zk/6NsVw4oC+EscLzgJqtd4gdFch3NiytOGWIL4zhHwDGN4AkvhOuey8pgTTgxZ0
m11dBkkWUT/hYUYN2T5vy2xEXlbzNoP2TBCEioch45PM5hIL9xco1ZARB3Xq+N/LcUXFAEOqwZ8L
X1vDdOdsJwV8HuZSNb7zVuAIU+i+Mi/Qr/4chKkqknRkrnr8wc3RaD7ym053MbihheJC5jqOGrZW
wDnNU5gRNNS9FrEar7n1vWDMZ2+pKStpjOfiqFFH4Fpa1eCmO0fzIpJBISRZbz85STZo+8tPZ1ha
vfqeKIJJPpSRoAPtFp4FDUa+cNFX1dVlJipj2caSQ8lFPMChZhbgs7f9blPgzfBzTQ7dUVL9dV7V
g0wi/s2bLPq3AJpiV5gwjv9+gwHbrek5zf+HqfZ95qVreUDiNmXa7wTZr2rsI3DVedgc9zushLWN
92HA5JjQApM506R0E6Jd/vb+pqRhbRdPhyB4k68gIxC95qXW1vtw7aDd4R2JFByF1j6ZfHIqy4p0
SKmD5ZBH8bgqGBiaEZLjHWiV7sIm2kywBKeRI71qOuYMUBkLf1fNcAY223U27GRkp2/QiE/gSMRz
Mw7oVcD5iffDWN5E2GMWuXd4nIMuBdv2Hq22HHPcO1X7pDj2O0bx/+4+VBM9fmTjAIpoBfbu6nuV
pg7sUxWF0KbjgiLtBTIQJvMGMwEmmKbmMgceUq30K5TCK0NFpWvlTp8YUA4T5Ge4FdNYiOLwiHHF
HRqICJ6sXzXi9TdPNDZBrvljpOJj2Gv76bB6qHYfJFNjQHRctc7/FuLHdUSzV6mw0Fdh4uizFAvH
LHzeIClMh2FZnLSMXWcgkIy6mbTLohSgJrfv2OFye4644km7ln2kXnHuLbuC+Sk1bJD9ZGSt+/rA
hme3BJPQRdI9ueIqm9YTmUBfBSI8pry2vpDpxw1Li7EqvgyJAiIL1SIIAuN99dhMoR82ukioQ4ki
7wBgSp2VhfYAtL27KKhNdUMYcdKuCJY9U+sIHk1lS5Yg4Jl3eUGpuOazDbCsjQm1Cvfj+hUkkAz4
mGQqiXDEk8720BGVlFOOv9qqFhW4G8YTz+zBVbZDpcw6BPOoicxBZYtqfLyOlo3FyZCBIMZ2zGYQ
EUZWs3EjnknEdC1A+4FFv6GGrzNUlvaGukWfOe0O4Re+51j63/73lodxfe7NDMRLP3DD2ixDRiNt
7tpC7nkb+ns+yfjDCfZ8Z2j5SoJ7Yj01FzevgRdAWDs7tp30nWnZFVqqHtdsxP0hmxqq6v16H8wI
THir0v3wJW3HBZBDaprfWJIoCKArwunfWu1M4vKg1SXNpOslMmY8FdihwqHPBgQw0VqXnNteYfHg
89EdaDuEnyEIqIym2ZhNnDf2lqTTbnqTRUw5mYkLWO0A8onlBr202qSAo69D2MIt+fGWRCbkjyDA
lheM7GsQt6ItAitgh71oZ86qL/NOgTY85pPUhTCUc2LMrDNBxgJJEZ5JvEG3cXloXtrbCQEzqV8K
1Azs5slMHtLnrw7o12n6mQHRWPfcwhcT6cZRUGZt6+zeLFLYGsr74wdMQeD+8TZEU5x1ozMbv6Ue
mZMmwRz9inw1XYDQVQcPnOmNqkGaYaGtGQr731qYYsxx/ODd5dpD9FgBLtCWKn2hjMhw9sMIgGAK
n3rH5cgKBRV9mqJRaspp5PohFIPbGz8xnwwkb4TYt+v5uvBy3hhRt1MFtsnMkIkdbcRcUHXfFfYV
LrwARNonqwcL3SHDKv3HfwSX/LsLaFN++atqfEfk/xAtFhxuiCfCG/qIYBgzpHvD955utJNVONhi
fqu3vmGGiZHloNTJ00YtsNsP9jAppmgJf7YfeX7UvC7iEFbcxCOFphUguSwJ37lIIEaBb/tmibAz
fL1Mpz3qJRRnfs+iQ7oCOj5rCYCuJjxRoIqbcOBB7zaOHDahjMOmfUg7ISKpBeNUio7uQq83afh9
YNz8Q1+H636cBbTwXz0zl+c1W9FtZHBBtSJ4G+6iO2czgb8JIP85jmC1i8pnaBCZJgeJMJpGPjIy
RrC78RcsdF18FkK/0ecIpRt707XSkfc/txaa6ije3fypS4S/s0GqrVwPsRWuu+NlDzjvLmUlaDwW
4J3tctQUcwzQSbIthrQL+L06skKpEwrQa/G0snCfNVrSTcx++8f7mcx90MvQZI5QBjMlxoLbkSWc
bT3K1odS/zHckNS+H2x5dGCnwDF/Ngkv9S68RyHT465b9n4G5I2EbL22Db9h7niBLBA7GJj9BqIO
kekFdTK/cegKJy7vNvJ01XJq8031XO6U3yoEYp3gdafGTXWLJqeCBgJNgnV4c4wLGe41nk08uCxv
XUrbm/plU9SdQliR4n0bILgJyY1wQXXfJ2+E8U+K6Pwe2K9wTdNYgqzHxVR3apeHed/M4Yv7OyxE
B4rZ0DcNFx5m/nyYFuIOqdieA3CntCzNXcjXyZOsvORMesK4b+g2b+dh8B0HZZnTEqdtwpw/C0qk
4TCaTwxM8ifhC4y6nBg02mnc3YI0LRmv2/ErTc8AbOfCT0sj+JcjL/ujrZ5+xJjfQzuUTC69HFrl
x+V85vtPzwpzgl3y6Zlxe+FmCTvmWl9FWP4GvquAJPWC6BjDa6shUP+E451iVFJPUN/ce7PSfISg
bcgokvAA/K9cRnmSDPZJxBGz50UGxLMv0wvmeHqNg08+jA7Kea5mlMjDb4Buuh+68LPJUme54WRq
Gj12RWgO/9KdtLDNeX1vrWyDxiutPKEFFbwDJKg5YGb4s7MhgTdgAN5dbUI1wgKxt8PLI1drnjB1
SM/Hc7+gdPA68m692WDnAo3d98NuRNmkt5ZRyL93xQ7TDvwtwgpk2zgEM8tOWiEsyBiw1Pbb3rdO
NOwRYkt7x2VgYsGnXvSQ3opnnTrCnEt7VM4NzZDvkg2GUEMpsTCysTG7fM2zWFKr1UHH5ZmJ4Dg/
gpZsIHTYzwmAuSt5lPFZ4Ym0EfevEB5vcobI564T1rmJ9+GdT/rLSdo//tVed685epuyobYkM8PB
wIJpD8Kr3YnS8fyog3gb6LCfBNziRRj0+NKDnGoEqecrwDm4g5NnGp3a3yAgc0f1cwCTKRUijrFR
l5Az9y/kd3arxHEbn15/HzmhxOe/PuGWdAus9BqlOkcbK2ZRPxFLCYBm6OSF7dFbs9XcVetIdet9
8Bh5R8qzGkr5KMKRgiu2OkeJ7bLFiaN+576z8n18rfZjNOqwzKU8Ic4RskhZWbwQqDKSbHurP/aX
ar6IEz8QNcUcCJ24fV9VoHWGBjMoeYq89olcgTlAKmY/VeVZtl3XFJrJ/aMRXHt6WGRpzEDS8Iih
HQqqvU4lPWxzn7igeesVQ+P+wuENx4SUmc//Gm077SKaJBMmEd8kcrx5dQU6DVXZ/yargOy/sqV/
1eYUadH9y977modbqEnGZWIICQsU/w2nWFlk4R5Stp31+/86Mee8kBpprCQuWgJS+Uf4Jhn5dbt0
NV/OVj3Fvybw6BIHtg7e8WN3/FIRZnstOmUWXpwN1d30zps5uxNCcTI4QMDt5GBccs2WNY31SSl6
3xraIEneCDxyLct4lx9EgVyoveNVus8G6fBFguMwqOeh138/lI49kdGJ2wfVb6hjCuQoV2f1XsCc
xFdnEzJCosJNAyUyJICXWlBCwpZPfWtuRuw8GUSBsjPFxwAE5cD5nglqiaf9bSsvHle4lUYUJUBZ
Uo4cIkngSLd17jH73xPBiSGFEJJ7YnFlAGZ8HZdXHgADsqyU7cAxKLkb5vjTRkUiX2I5XUPHyN16
nZCCrjdFPaIwm0dFcURipX4DUFGnlD1qcIqxBPg8AQefXcXWll6hg+wfoJDtRlswfEKr07K6xCQi
OREcBO5mf4JFhtVy45S6c0/rwafKS2qLhgMOPE8i0PH/+jEnEeFxT6kMXzUJFPoSeLsqHYfcZGR5
vFTX6iZoDKc87M5GHZTDg2tIqZq9nR43ONlnEYF0IoVw74WLcTN7TbT8XKZmSA2s4Dk17qIP5OkU
OrM7odQrWefWMtg7tafzQSzDtRJ0vqJWNDzHCyJG7KO9IL7t+Km4LPut3qTAM6zur02KXQsLQrF5
5Y5bv+q2yx0mWEZ4P0hsgIRgj5hxsPpza8r693IvyoZ53Tk1YIl8tnkIMpCkJ4hg4yg0nFTGyqid
E8CffPElvm37LHtbCQfoPEZFiuO7jdAHlSZdQsQsnb3ARO1UPqNQr/120dG+BTHZofgBEHiS7dqO
PPV5csOw0HeUmO4voPOBZIDTUb25worpaJAlh4HCVbkXPF1NR9y0fwvDsZtqO6ijwKYxj87938wN
BKueokBDE8LSY9IYm9EUw4/IjruoeWv+lpUqs3FFUuOejcEWsKBmIXOchfEQPHMdAOtS/UnAQvbC
089WPZMjPaYk5eI53D/WOOeoGxYnjrVJEnVyo9n1QD5dU/U/oGzhXCR9BJZttgahzn65EnI9eYmt
6QDQ+cGqS+3/hrG/LIRyfvySiDvD0uBO9lcUUmaZ1uwoi9C+J2YQ2z4vrLeujT0xGfr/yUEVyuu9
gaIjZz+ykI7/tkay4MNaNnCFL5M6wxbbBiA8f2WWNqlnBixz8HGAFJ5QgrVIf8+r0nTwcim+KdWU
lKO4wPnwbF3L4L3GzXkT9H1lJL8KokuVsgGP2iFX64q2a4QmGs0+31nIacrkgeboKTD6OAlmJTn5
jHzC9Tvb2LHwgU2g+95jXcTE/2+w8q9KLIMo1mHxjO8wAW29T+z6ssJzRdGbtHk0nMYVzC0KIjdM
jNV97EkvoNMKiY3OCps7S534WbiUSpdOnNAPJFUf3581QEmUjKTBJEjia2ZOD5g+11qboqD0YPsE
WOQvTXxUEMVogd2NgqNM++339u47hnYbZMBVgAaMXErmkDca/xbeWayKxaVs73+Cn/r8zlBZLJJa
HLeNLNCeEUE4x01G+HLKwPC8YLcUHUEjzaeZaHQ7VNIe3sPezVYhHgiJ/mSE6eYBSUWrLVuALrN5
0e9o4rvxx9aZgrvbwrQW+If/1ThicA0cPNhn2FxKhNzI57nhIyDZlkv+DrEHgvjeQrl2F2Gw5Gvs
i8nuCYh0BX7ZpH6JRJqBtBduCjR4tMcjKtuY0f4A5v2bpCOevbnUjp7et4oCE4kIbWmqCd+RN/s9
J0aTIWZLzPJelSX1sgWW7FNZdgPhsCv1M9oQrN8Bbw00pJznqf/kGMO3kXArz+M3e4XLcQIZXY6M
XIeTJ5Q7lHK3ijh1E1uvFj/G19E2ES9a3NVTW1iiGhNvXzflNE5J4zzd3DvuaepmTp2jUoU5ByRe
CY1jeRALGiRDJWweH2l1vacp2sv4MpAo5ZVZR2IzboDVsJoFnld/nON1sOrtCZs+gYiHI2Mb3U9j
OOBhi9qrlp6irtMzi4uGlzYXe1t6hRHIgew4+fgr8Q04aKOVC8dF+Kn9IkXGv5Gl4ViuAgNsxSyt
TwSlrpwXZxk42lCnMuWE74Y5FWtW/QMu9zFFzQLdQnd2nCQNgZ3tqupblztfJ08YUE7PHGYYSzUW
h/zhd/+w9cnsqDqz+e4q/LjVQs1vU/y3OtiUxpRXS4QiPPduhaqtHN0CpwgthsRq2VdSwXjtFRZr
S65MOZgS3+vXqnsu87Cfcxnd0MPEipt/dFLUNc1x91iiDOaZwwjp1iCuvQ1RpAcngB/RgasA+xzx
+MakMLUKoIH80wNlR1lC7Ceok9Nxmsblz7EvDQN8c6w3LIQrwufEFjvZNlkZVljH6dDl3wWNVwxp
mf6X5Ltp0SrhDpZD9aFMEHC63ppbvRrSicIdXXlyuzKNipwU1r+Ed/8BkyAXt2pk5VJ8TiOJoonI
dc4qjCFutK4V/lR42QlQfCrk7XSVk62hwWfpyihxdqWbLmf/Ok2RcY5BOsACBALINv6gcrKQpfZX
6IxTnnMOHHlh5PqwvL2kEXSBLBA6nPI/lrALxpILtSPn5gejABFOF6BXrLih6yQsl2eA64SDRnFB
aFRZnEpjqXlDE2z3AZ0ccHHM/okfUzs9Nqr97T9g8bReUFV/YJqRMY1RwjmSh0C43+B0eUD4cl+g
HqJ+bp8CuY4RLjkHSyRpOzwta7B5CR6ve7AFn52FtOkkIcoGe8uEfKGbIfUOFMKBsJaaWqF4eMSx
mlgXUdXpclRaMZuq3okLj1r4ds92HiO+9DAuELV5AjX5T9lVjIFAbNx+uPBMFElyXonyNii4uWFy
YYWgv/joldj3OLcTfDnjc4/NDBplBdH0AqzdjjhnfEi51trLnl6MrUvVciCSJ2sGUDvCvwK439D7
YREYAhc2DL/eQWKC8XsTBVWkPf9TNplefTxzgywSG6sPrs0KYuMI3QxMv0RsnMNd/ELp1teASiDI
wY08V92ycPEN1L+tBpaEF8ZGF33b/ga7MHmTsCaE9QacpHgSCza2CumEJHL/YAWpphozpqEFNCSa
OFICpr0/EPI36AIbZkemdm2aQRALAu8PzGS/iir0nMpaZEc8VTwObMvggRzNlNJZFlDPNLYKJ3oZ
dKFAlRsTpe98ZDpF8hNaWpoCCYKe7m0d1wHdugv+1jE61utZEQesyVs20f1n6yd2N69HlSVAgfc3
YMAJ+k2eNb6k6E2ZssTNLXK2BSP/DpE1YW4H86x1ohd83NciwLmY71V0DCwJmDF8ym0uQ6gAShDN
Beeqg9CErVEpHJDpEsMKTRHL05D+551lL2PjeAtpnmOejotoC76T4NbQHkBVJVV+MCHlwn4SqPSL
ebddvwtieuP6focpXhGgmzpLfLrQzKbalZGJTjbIAfbpKhghGENACdOu6fhvH74rqB1xaMj93jm6
JRRk5jZMZGAaJeGPqEK+7rX1U+pDPt5SYzhl0xR5y1bDag6FlSDWgDLXeQTZ9g4LlsdOrgH5ZdEl
THuXfCBkZ2fcxmiLWlL1cK3JF31KUZKDN8pV5Pn+GMdM7uDEDK65xZNyw2LJMdCgXnm/bwUyjrxq
fV5+BFsv2sryg4nLOSaMlRbfnrA5isuNPGyeTyixl3JmvSOHettNtncZPGOH5HbaSBNFpMj5Swzq
JC6TzMXACB51BJQf+iYQOQvXleM98JyggfCXNwqc2zlfF9gNegainJCZZ73ei/pqaIX1Lf2o2kPx
0F4GWWTr+gyb5ZxlQUJoGtDnuTnBx8GO5sEeRimxnKLWEmvZqtJ8NI8QPC5X8uLKzMYGdL25BuQ5
7RxWXvonVX2EL0Z26orwbQLSzoh9OANbOxtk03DAkhY/ZBA/1x4wMSi9caePT4vXarlHhtZhNXF0
RcpZDVjaHIdTYYoEGLInr/qiITU2Uq+cFLdtlrm0+TiS8QNZjjnppwVVsK62ZvKeeU+kZ7euVjwC
E3TfUJYvqIljPFOiZ4/FxunqyeCRE1RKlyxQu9QdYd+FfFibC+TbybwSnggSYngsQTPV+YdwrLn5
LVxJ2OeMADR6UKCXDoCYw0kUFavejlhl9JMiqvZnwxPeHPF7gjyQVRW9/z6Wn05IVxNgNyy6UvGp
5f4zGGHShddMAq1Wvg003XcFMlhKGBMNTLLCDTqAA5fdLmCRHJK+QXmj9vrWYQBypH8DEOmU9P2f
ZBUAXnsK4hi+8hQ5wnAS3sAp5nQ9lbjQ7jqB1yifPLCiVMREzfIAWXyYtARKkuHhQ+OrVGvWlBG9
Xq7uTK3QW2b5u084V+C44KxJNKYmB0cblaCLdQP8u8Lj20N6bGqkkJ+yxYhtvpR3wG0jJsa7zXVP
n0Dk0PRwoD4TbeO0XDTctXK1K8noG18QTnPgzEeI/sCGgNWQy7X8DGXHawVxNcvMvHMwf8n/9+5o
SOAW96gMoJAow1CqlQAmMPgKZoz++tJ9IjvxkQ9TQWgVhAy7RGggy8lOCx+3tpOHH70w2xtnCkpR
lvMsYkJYVn+U4ora21q/FTTLhSuZd+ttNITrLP9F239UItbJQkEB2+y+N++vpQa9DSrVRUQ/ErJu
+PVDGGAcQma4SxcMelGp8KV9ljaet46FZts+HwvPJtEPOm+Pe94gfxq/3ZNaikaW7/BUwPfJGpMK
gjOfIcASJM6dR8uqHGTLvrsSLbFBfXdv6MYY4vPYEGyPbz7A00XvZsrGhk9l2poW881gwOTEZbPH
vg4dAXc15wHo89K1jgjBNvH3auyAElKy5JW4y6IEcU7+0ZXHa90h2MBl7LdhJ4kAofv2qtJcNMPE
YVxWIJvnylyD+baUNj9eanqdFuuy+G+DEP/DntploKWUTTYInJ0TuuFx/0yG6yOomgYt6ZXigs/i
4r9PA4Ij/FqDd3PvNYLXNzR8373+ndNrVtVEsGle/WNfWGiXBcnrRupefivrHAVQIUUXnvNa1i8N
pAMB9k+K6hrp2hVgBVbGbKJn2ReeIO1wrywaF91qA0mRD0E8weHw9HOGnsR2K49zLTB11I1h3Hn8
Os1HMPFkXh5wlyUzJu82Vml+4t0NjWB+eBRBP3VtE+JIQBOVOhCrUudQgNwQY7YuPZUDXafhZRq5
FZgTY66EmZJfM356BsUAn0MgseRzKx1XvtWCBKQ6xvu7mEcLkFzz0XZCykuggnEeojhnhHsVAsAy
oJlkBcEnOFPagH2QcbU7EHZuvDCxQuU5U5QTPNqByGBfQNJ3xeSuZQ+E4YlyX8jzuwYE8jsA4UDn
L579PzTvmnkRPlmDwwxUOeV/awDuk4D6UUK+XqD7yunymuakgZeuEMdezIa5WsOakpwfpwXywuzF
UW2O9Pe9bUENXf/s7xkK+CarVaO0SKxt2SNte1uryeoD6uYSSxKt7jLbMX/OgRdM385YxxkCylaC
KJ65G7XPAYHG3fojHuw/4UkumjghdGt5V0V95rxlypYFrc7zIm83YAoPkk5NZgYU9hatux8SWUKw
JNEAeN6gsRlZRcsSUZxPEkrUEbBUdWb3yJGJEvjjGCjWUB84epVczFslK4kBvTao86sqH42ecnZE
vZbXgAIYorWiT8B2K5wv0/kV2jC2Q3DUlk1w9oOxh4Mv9stY1BYFe/2ACklru7Umt+x3QVNyVfR5
rnhc7W7gbV3afa04ZmxIXGo2Xyj4tjoK8hoaTEhraFNZrMpKk4PJEsCZHLytnH/YD7TsHqs/hdUk
3RzWw7UwyzjKCe7oBKW7Osa0Ea8IOJYrn6CInV85ShGia6XeKGOxc/UHvPUusmCAWhGAuxBU5ZLO
QvWYvueKS2h6zxYz83KlJpcNGoEvgmjSSqLK77mAQwGBcf5MjaOpWDlhCi8adAR/gLAh1SICdYLL
Kfi6dpqEzkFKSXslVFDyOeOSAjfKLV9uG9M84EMQKedq4bBXehc6sm100o20gLNPBM6dH9lJ5gXP
FOS9qyeskMlxZ9iWhTJYjM8cNEfIkslGoAw6f47js81kyCaHNxr0VYCgwAKEvrws00GHIDi8S4Yz
aQ0ZgAUUP0XgS1CM11LgZ60QCcs8lx/8sM+zFukZG4VOsj1p/jgDdEJpQyG3tcX3kkVhYiYJ3jYy
UbX484tnyxggPow6/ysAbzZCZmLdENWI22rESEAin6utQCXtUxF1CQrpsYWDEJaIDn++bSJuB6rS
zgMtZ1w2kOu3sX66rxIg9MQyQs/MdFdTgpZ28a1Zys9nkRwBoGae1W5sWoU3PWxlRlUUUN2xinqr
r1MnNJZjmBs3KzU5FvHmuRRztoiaytxHR5n076GFxDBxgZy3xpyL1FzGaL5PGp0QJvbQAVr6AHQY
eYVPB8ulO8sQWEX8iwU7FI8xQktad3Q/VI7yOjAG+wNCRx75hW6OyHalYxtfW9gzZJQGidSPxAbH
26JoVEst73He7X1IyYsdJgm3G7QQRx/hKr9OgPpY5IGV4P7ZoXFKo+lp/NQPqAtBmNJFhQi27bs+
JgL506PLNm4mBy5s2Y4wvzw3Tzxlo2V7baot7Mk2gDAGS34OszS7tR5kU/87crNJvB3kx6ecIv7A
XZL/P32Wu8FcXNEeN3Z1uFUWrtFLzV7l/SW3PdQx768uwNhlXVQPE/34yY7+t40V/O2Q9/sUtGv+
EQNVyzZH2Yl1Oy55dzy+uiQm3ESVSfPZ4SJF+Sy4ROOGU5KWKo0QHcrh69PgP7llhs0nuHYAn4Sm
EFa2SQfZCfp6x+bAbsQSPzw8okpYThY104YrjGg4GIxKEh7NEEJ2STQ0wxP/Wn6D7ZIoXNs+EycF
TeBXtLUufI9JUETJ7XKyuuYIkmg65gbRDz0E+SV0l2Lz2aJZ98IxbqTkR4kYyh12CTgRgxD0+z6+
762D9Mj7Bl+lCT0E88w5qjDCdy+MXOjIfAL2T0mUfMN4drRE3ptNAAz/yYUEAvLYpk/EzsK3RKm+
oNSNhE6WRotwlghPk0szvNwcdqkqKtBC1ltq81iskCG/GFA2R5WHefvP2wCMGLkniQ28D6L0cnG1
iuowNvw+u9YcmVpHyYjSHIctLfAkelzwDW19ihpXOXoKXtdLd9Lt3YlRWMpADxAI6wr2H09jVmys
PsKjfMseAKGqQmCTqLr7x2D8gmlrKx/SV3soq7M5tozek6tcbItOw0aZ4tZvdZalisQrWFnghz/t
UDTlkuf2KfBWALCRGMOoo+hvTggM+VjCxGtXxxpc8tI53Z94RMfzpXkJ5X5590adadMtTbnH7ok+
n2YVSdih11mryi6LZ9VXOhxG15HEPLJUzwv/nZlWmlmEczrpc+bXZGbbU0wXu9CAE40Zy8UtQaIL
mOjy4MaqLOG2dMboI6ClEufn2dn9BbH9BxKoyoVbF6SVFp4P8rb3RzYKrp9GPvtOxpra1NeMUZ/V
BpRujz3wRMgbgNZeDUSTNRBCD/s1pDUcL+eVMYqK6FV7ja+6ktKCmk/tQWvieB6MNhNlwicDeYag
E2cPmaeHqVkMx1tve6nB7lEI40EGSQj3qTF5BHzjkq6FEv9YElgHzQkHyIDuMFSWJSxqBRLlMmg1
uWBgrASKOmosQnFjL2tQ8POY8BXTbD0GlkYJY4HoJUNtF5QzC+FMxP7pmYt6iONkpx3Uc3+Fq6YC
cv3GbtG5hyjY1mViWB5qAbOZOx+NHqTeM2sDw/8AQviSp7NrgfU0G0584ewoxn9DPyl46IMxHoF1
lfD2Ov9AMOizSyvIkG7VkXBUEtVL9FOHOUGFe1RCxC30f9pUGvDpl5rCjUTfltcC7HctpKu6A7tr
d/p/PdiSAI7vmtSEgbJK/TMRYVx/FGFYLpZ0WlS68jZsnrbXnzrCM7XuN6WjfY5BesOIB8xL1o47
gJLx4CoNI99wN/m5xa2GFMtXZwZWTiIkxigL0b/hn1JklbN9bKQGPhOICKlABAqghSa5uwa48qV9
tvqC28zCO9sdQ4wspa0/tCYbJRw4gp3SloSuO5JgjB7t+nW4QeqOlNidhLpu8Gep6wnxLJE29zxI
dqKnbu7jSaTtXeB4QxiZNEIul55Z2DenHbhnZFtsHghn8PMo4c5c1HUQ5KFnCaHSAhPjFbUniPlI
HqtdVvJO4Fc6nSStF7TQUCK9vWDuM0wjKnB82AzCh9l9qOBgHBr0K2GaRtwDyvrNGpl548gd99ey
y9tP5Gon8uirEN23iw38K9Nh8PTjzdUrPvd1hRh7oxqS40n9p18EeFwVxcaTWu/D9CYEGqxCPOtq
7gS01tO4yqyrk7XiTxn1KjLmTnRB6JhlTj9MAu+6MjD9oXsququRlo0JvW3ccbQKQedteaZX4PTy
FxCcjWOulS2MXpN9TYwFSZACXF8VUjE592G0RV3RnwTHhEheZhRw6oFzo/Hfb9ueuePOnIG8XPTT
g8IlLQGlHfXbaiQ9b7nGpVoowt58tJaDnl7yC6Zs4LCQYLD8t+jpncRwWg8drgjUGfKO1Dc6IXxS
V4bF73cCN8x+FIj/3Vqnw3tG89aLMBYxdWNIprYEP/9f5wd74Fa1XjJDkPY9D5jhE+1E+3tUpmvo
cNaM/xInGS3uSJf/hYFNg2gmWQphlO2uF540nv5fhHWP+OpkVG6OicN4Z/umiPlMjeK1wlNGHvfj
BuwMa/+IBerxh8OQQg9wfmZns/FLQLMnI9eW1U04bP281po3GHLNAjCQhv6LPzd1JvKM15+4+PE0
axMDiM5dlFcMY5z98oxLfH/EQ6932NbyVNq0YyTZRMbi9bQe2t5ql+S72Cu5LO1Km6gzYkKHARLQ
scD20ja/rJGDqE9vrTkokW0c2X5v61NktkspAW2jFZIxophO3JlpQ3rad6hbCUFCzP1QPrYnNCcD
9HSmvDzytwtEOCZedb29knmhm/5sn53K2zxB74bn2yWlCQlc+MsaKbTA0XLNYXd9Jb9BgZM/d88C
d1VWCa72aS/anhlJNoeckeO6NX59CzqRNzuigcP/GuE8u/8Rw/huP9nehyrkMZTHBtl5I+1HUczH
L3JliEVFmbNj1E89LGIKnySFxxY0tKyk8TkJVqJn8juXb4WOuQFNL6Xzp2kqmIYoWzH6uho5WHyf
/wlDr5VSlxaM6fehFhvFBGi6gR/V2HW1jTUB5J1hpviSygO3XQ0Wp00TRh4u9T7m5/aDsWna65Od
iwVYne57XLYljzWFvNgY8cwpT8Ih6Cdla+1Jnn1HLKOzzzoMToaTrmT8rYmcy7mgaOMBG2OZss9K
GIwkicmhyTHVqPT9iUUsXb9LAl6vYgvMIFi4I9gwemcHTtR4WPQnXSLcPOeyPFV44sD1K1WOOhnA
0hLLUZwNAdEQFH7mj3QerNad31jQcR4GgNtNJ3kMk2amIzkSHbcrbV9s6akz3cKmDpYeCTS6ZahE
cbb3Djfey166hkfjrdRSrViZn1pQBSAuJaU6pe0cf1fJ3JlVKeOrSpD5GzJZVgCqwmGsE92kNHGN
frCUwAjB+YwkYPZYcsKuyujMUZ3YDCBI+EcKdX0gKdf1k3n3rYv8rSs+t1AOZr1KURp1JHZKBBsQ
UYvHBwqmmcWvwPwJQcKNRFv94BUIf2hJlLfnMfLTPE3ACDDxDneKBSVXDAl7F/fEAcQMJuSjXakd
y8OHNSTQXyUc+vC2OmrjMPnrPKlva38icFhbOJt8akKvOwpeIKznZB3fDVuPCIfEZ0BkE4DdjqJB
XBrnrmIUe5cc3eTGc0x/wBYI5MNmrUh0QTlVqd8r802W56jsqqg3neP7CmCInKorYkoQH0n75mb+
XetknATZt94Gz3TvZLwOXaM7W8gZsqPX0z8jRELkdCDK9PEPKcqD+vfSj4j8r//UGcnqX+zSwpyQ
/u4S7sQYPSZki8wslmyBjXpkSajv5BcP97MykKreAzf9KGGVPU2koODPexwH4Km+O/+LhhQvnR2d
JBpvdCTcszgR0cJOE7OGRHiN9ud/JeksQ8Tty4EngG7/AKMxoN84VzP6fdfYMK9AfHydxllxrz0M
TJ3fXzbKl70QvkqlCXZ00K7gAfDPSTwwGrHpZslBsWqdiXMkW2Sm+UgOeop3VrkpUc+C7RnnRkDK
Ar8/WkQgW+RDVsu2NdO7JkXLmwMtItegk0tzPZGSasCU/wspi+TsvyzJWF2roHA5QEZeWx7BCCUV
hqBR1v5Io1+AqSF1GrHeq6ocRHs3SJwAudpShTVyG4eH1vPBRKYWY83PMGqj9wznWJSS4F8FOfJw
FtJ6Oiz8Vheo088vSRdyV5dr0zgwAX1BS/tP/PFVfv64G+AZ3rnjeB9QLxK1Z8vOn/MAhEDP7Dp/
QbxjeIhvYvWQp9Ac9lgo1RTUx/rrMZiMHlM4NTnngPW5fEA/hSghh+dYxTgTn+xqwKGS6ChjO5Oc
lxwaIngU4TJ1i8JaNKlPEhHPP666RLOu/RpXvUz85YWWtFp4vURPfGPtJMChFoB8JdGMltOafBlM
IaM/MPntXBobWlxanTDYiK+FLkJ4LT8STOYw9Bi2XwWmClxUzPnTuPjSGFBxzz7bbMWwROu4NTTz
AJBkMXrHfSz7Dv5lYBHXKnhzM5l2AvfYB+ag8GMaQfnO61UcSz+CDeIxTmZiRYtP3OoJ30axyMMg
z4vtNR4dUrydrva/PznydYQ6JGmwlp3OMm/zknSQGcfQ+aMU3BM7bRcZkqI/rPeE8krME6FXDQfg
EDRc/kAzxQ8v78pqlZVd7cVq0qF5gi0xv9OpcjYBh6EbtL4/wD2vyKV5rRrZOVB/IuCWTco0Mn/f
0itE9kZSdnHkFEhEwqGDllafkJaB/14lybtGiGCXrjyL14GIi61wkyQq79gZ13eHKEtrmxsFVO3+
PoENFOUAyoWfPWifUmefpMvW9SrBrUg2yZtRQX7Vne+BKmD2StfPy0d5MQJe/wZaz5slqKhx5H/W
vJvGn9qu3VpY14wjlRPg3L54irbm57yoSBi0/4MoVN74Uhjti36psZbfSF1+6rjTury8SwPDyodZ
p4c9gFirQ82xNw3ADmDzmjwrOEvgglxpUYJ/A1Y/dz0aOR9jREOX+0hAqUAYA/zEWZyOsAK4xkpt
M+ZCt11D8cJkRgwZ0e3+N1T4OKYz0xeiWo7/9SSc4O5mxiGMd5GW0cy5Nhao+y4OtcakYzGIVDsu
DXtBwJGr1l5QImJpe7Ai3wxJ/La2ZiyyLO600dO7/MMfzc8PxVzBNXQwrPiMPuetp0EZzbJSPTo+
1am51KuGcw8vk4HwTnYnO36UYziIz/iD5phrrQT0xRogRAQlbHKL0CllmQZ8E9dCj6J9+7A0l4Vb
dxYfzgn+yV/Pu/ajK8b5WT2b3oK1RyCsf0Af02iMNs0fdinQDb6l2zstkCNtzeGSC+1LRr0INaNc
ADjN+d8/VAAujdomanbmSNKPk9yrZ7A0OvhWGCz14FTbxwsQdc06qVMygdNWR4MKtD0F3NHcmkqs
LrRmT9QbNyU+4SM8U3X7r/rBnLAAU+jfiuGYMvKSFYCJJsR0xfHBCf3Iu9q1dLGcQnLbeOd81vFT
bWojsNUGJnygzoRIiUXPcGpmWRTtBAPZtQEa9scilzytG1WVYZBc1KPgOWVj3pLqSQmlLXuBfdJ3
iVNqlOP4BXSDhBvtRgOa59ESxQ1Ketvmvk8Q/B3i4vaqB+TRDgnFDPN4egG9EFR2aOI1q1+HaIKK
RgLdYFb3D2+RJAQI2vrOcVGPO0JvpMGK1Ms0MZjIHiifcfy64MOxAm/GD4GO8UrtNiEot6n6mRAX
Om0wsYQWrlEnhGDs+cSexYqyCbX+B+XRGcuGfQh2FWt0bgRmnsrmDaG+DCijYpzvWFGLhdB149S4
glWgE8E0okZMrT9w1uly8natOkh6WA5j2K6//Q1V7iMhtFVAiO/51L0dPA5oExOfCz0JW82AwT/Q
SySC0BOzNVSrqLtCMc0sT6Smx5iDdZ7SFkco69GQAkzpf5RWZd3j4Sr4tq7F2DkrZEooHnyfHouJ
JadtrAgVCswsm0AZsa2newoAzTYeKJkbRQ3uNqi240Hft8pLJMMKsiHDOp7+Z11OAuAX+WKPQwsg
n+fHiS5Rl/sjw/ApP/tSJ43xHMFlzjdARr7bpfr6LSipUcmwHQkPxgMTOLl5EjvkxkYmz9Ubt6sX
Aj1SRRDrK/SZTnYm7CvL6fRluCSJVMIe/MKSs6DzYV4BG/SvE+OUF00EIh1jcY8NjrNFwGuPh1XW
mWtX+qEwZxhMOCCcWA4I8fd/QoroGNohmZuQdTubAJP02gKzzf9IOtETMQta5e9fQXIBCASLeG0g
49kJKgtCOBj7wsCR+iRpEV9KkNIpzoLoQeZyeCHHx1t19ijmvd3uxC+CrcPmWSWQXdsIRyEIwNBD
7otmoAvHJWgJxdFd7rOhmVwjkVwwu6/SvwbBKB+eDVpalbB9fZnAOhG07LgDsTFZbdr8R3sObwC0
hXyoxGHpX+urh4xhjyDux73B66zLBxU1MOqlx39sH8REz6rMu7p4U6p6x+XRemN2NC43gLe0/Grt
xEq1mR9Im0omPrcl2hUykoyNe5Z38ihlZgEmbSbh2eiUt4e9S2pXJmTSfkuLrFOdJudXuHoyOH8K
6thdJLX5N1DaQp9xfAGu7FpjTs6B/8zM8p/6o80+V0vc54ch/tvsaXJj8esGaKbFmJQbxTSBPxiE
A/T2Uk7q5ow7tHVupMQ/9m1K3Kpy8tRRdBetmr18zUKKW80urbTxXfQoVZzhdEGJ/j/aDYopwLv2
3a9VhKOpers3dGFXcPSpRjFWJdCJcX4inALdz/5LtdoKgr/vab0BQP0hcbGFB9TKrxAmpoiXDZv/
dMa4pJEI1n/Lb1xZQHmf8L6Zau8lggJ4UkX7oLIJrKnIw0TmA5mSKzt7VSb/2VfipUwlXc+ZSbWS
B8oN//4N050pYwsKkEEizEQtykC0p0xGh+Svgy8PNaKfe5E13bnyxo+6/ZBsGOiWnqsVHOr4YXYm
nL/DRQYqDV4rNH7v79gxFUS5F1N1fI2xOtIj6r47RYlAOP95aiwEu2yKCo8cRmoudqnzrEj85Py0
oqXc8Zyr6+OL4nHB7KouUx6QcDuWzwsWro+ySiVgXEl4JaKmcfKFJFYTinKJonXYFrIOrlsn3d83
d3Nn3GDrzLb4ni6/fBNGu4E47Afy4slB2w0Q6h8nVtMxPqi3ZKzWLxGiy/34iggEhvlTOyvEhFuv
kGDfFICSZAFVf16zy4EGkRuH1ogDucfAJKWm6OMynCRjxgqBS7DKa7ar3Wtq1dHHSc1OyxPvRAhK
Z8J9zLWv12WtI17Ys5LFmu5r6lpExteim82QG2xlQ2QHWTRj8kMFw/KZnSERiUKWl6HwdJpVacaE
RR0tfvdFegbQ2o/+ibBgq3VYxR6cy9PXuvxaLWUovawtq8fezY3H5LXmAATauhPwN4C6hiUCVXe3
tr6GRQwAO3vduzxQVaJk0fIJvNmoLGEOhuvN2b0nGJpoT4zHVilLOxQNC9pFiRppchIw+dIK3Rn0
9jEzRySQVqLOZJzgV7Cq2uwP46ON9qb4nD8xYfM7mqtrQKIXYGIO2nTNaiH90QnUdrpgUtZ02/8n
OR4c4+36v4hGWSGdDbUhkAcErWEE1pForuOrZV8RO/HLtYMII9hRBJ34eU5jO7trdARIi5XvISRp
5kD3KgDjT1gYXKHt8HT8qmOhURAody3Y4oeVuPoxmvEnPzcGCTthvTEREzp9G+7R42Dj0ftYOOqd
J6vmuO8netQh6kAVU7g4dYMCqaOMrcc70A5uOKUZhqaikgaYLFZ4oLvnx381h+sTU6cTinaS90WW
sOqbXknM5dRED6dcia8oYSIX8SxFbjDgdguOD5Qu/T//cpXx+xJe38kEPvnwMr7OQ+0iwp46uptg
zuO8QzrsjalEc3f3Fbmzjhsdhi3FYuDv2FwdXyk0OyV5NQerlt3gmGPKREo53kkqp1JhwPM4As2s
iODvK3l2/H3pJPb+zaD51WkcfUp9L1BmuOc29WHH+1HZttRVSAD7sw8XVS1RpBi4b8ZBNNTecZ8b
2JzqMlpqQ09lzFeWS0rL4NAFFikXp0txYo+ES/SdLkcAkpqDZDrfDg3FcDA9Wuq9WO3asVmI45NG
G32QKLNjyTsMobBZtZ0QlD87pmb+ve6xBMy/REgQUvFrsxcBwhvSQcqGUvXgcNJwEg7uS4sLpTQm
kUki/Li1iEWQXD6lNYS60qYX3i+AMgRwCSv1ChnMHWkvQiUg4XxYV31vX7XG37hy7nX6jCMmn4q2
2VNTzkIw3nNz+bCTVU9f8wpuJsKDPWVXNVTHxusnAC3fVlo+/rGT/TFOufehgD/NKFUKNS3Btnug
kkRmzCeFLCmSsp9qGUqTHG8Rs7d6W5+gyFtK77ikvvIvL+dXbo3UzM9Ufd5GFj4uOAlbpg63NiTi
XR823YxiOh0qSwX6h2b4Tbu5RXYCXEE3lszs5rKY6uZF+R1yH1T/jx1ZYGsb4ipgg+UpIrXYttyR
nl2xtTndNqTwk1H7aKB5mc8IBjXA1YtLV5cgdp0YaaoKy3fNZOYzaexVfh155ahst4urvNUHfGyE
nQeMSdm2ZMqhWhai0kiT4MtBGcrZZ01oyccZLeGYVJrB4wMk3VByXL2wtwsIDhcnT1znzQJc7hpM
5k0A2BOOzkCC0cBYQsF1H/RLrFFL48HeBcL5bzTLculPFQvz+pRMVuRZu+TbR4g96nD1Xn0M1/je
ZTBaKS/q8zwmywr6FYZkjZ3nL6gvKJr+zmRBKliXFtV4tt6MIW2Zqf6A9b7LFWHrMSwDo7pKyYaa
FMxZQY9hnwq59ueBLJQcWYNEoPwLMyb3BiiHEReKlqFU9ERS+fijuV6GSlSvw3famxWWNyXj+YeI
86LwIJN4gPZDpUCNCC/J3yiMO/Ii7CUn3B4e0nWbdLJwaijOXkzIWMyUKSNiTwm7czqapg4gCKJi
NrguFcPMfO4VTMN7ltBLTmpwKdyUvkK5NwqeRbp45TK6axS/2L5fXsH8ML1YaY3+l+8OUjxEDlVZ
Xrx/7xUWaFIig4bg5VwAKQd62tjPVpSCfMG/bUa5Vups4glbEeC69fA8+CA3DFPpJbyvSOpNJ7fm
VxwM5xP0WbNtALxG4M2xWX8y0yZdMNEWig/H9alXygNcQnu691kCXex60FghHS562oaJoJ9Yo1QP
y9XeLB7hmFwGRYzPBYdXiRKNoFVb/Z42WffiQM4M+OY2vw59fQEp07TaG5L8t1brV28VQVTMdcC2
NU8q8Yrv7YXTOKWRHOaYIicX80sL63ax7Dj0s5e2URhs6WUQVxUtz68K8zyF5U4u18T57nNHw6ip
JQpp0GkGfCfiEENghWt7CU+v24QfhNqe7cKvP6Ix54t2HwLFfLAGcnHpQUrb7uu4cEuqpdtkDVL2
zWn9ouW7Pt9/9rO1YjZy6f8JhQqu+zZ4NlpGi846O9XbbsWTEjsApAiyh+plfRFbdn65akKMbeki
Y2SG+10ro3CdpG/PAMy/jNWRWmu5+En+k0EmAXdxUi/WI3+xVLxv3LVWTBwLHkTTcqIDb/xkBEs7
UwzDBNdjgW6ESXIn8BSQ1zvMfGVff/Gxrd0TPoVxFgD08MB4ydwIVnXUhkSxHfP0Wuob6Pn0r65x
ceF+Zq2zANdQqtP9JUyf0CfUhBOwPtMs39fBTie8jLbDo79wOJRKApOwrn8ej+4UmCT81HbfJVmt
m/dINZn91Z1UmqnvxLYbMIqIbb8eo0p/tWiWpmXre3/TWk8aCqUSa6Inn0xHlx4MiJQPtzLERdW0
9YPUoLwasjleRISBn56nEZXTXhq2oSU2I1jlWS2tRMAMtHajAQ7gXmcXcKVP1PYkgdTFfP4ILcoB
YYK9k+6iF5J75nSB0vm8ReR2rUCOMXAj+EgRp12ys1jbRM9ThnXP/3CkM37S3ZBAU0ETkG50fzpl
7/yj8t288ylY8eu1PJa+4Q62hQ+kyr1I8NXiWl2gEsTz0xRMv3py6WDDyiQG7IxnlRPV1+hQO2vp
6kuRBHYNIESiZ63G6gn0GBxQoKN9n8OldIAFgrlStb6b9SjegZe8K21tAzz2XqBcqluZSobD68RW
5stjlBK/yolUyNhhruxrQvJ22ZTp0kTpTQR6g0wRfYMaiQx6xqKWT+VJphAlMwi6aEIlTWJeSKH2
1n3PnNwtsJQMlmumFiIvhvEuy2/BlDooPN9rPf/D7aCKe3uVaLKTa/3Ps9v0w+QcxipY0DWckXvw
LGgDjE/Un8sLF3+luOJ5xsogF9rMCuEgHtM2NQQAT3qQksYLS9lxVKcORTDDzKnA7GaYYTzjYBk0
uPKlAVyMANQeK9n2/mM2+Xbqk/ZoDW2ORWp4NLG1oBBlA8vFYz26qq+Vp9SM7cdHcV6o9fpwCeME
DpyHOEYsrysq4p2OoQORzB1eSYw3sh9/CW5oQYLA6DeDVWz0JpYT7tPEz7ynvCwqHmpUYWFI1l8h
vup5/hlN6nexIbWhNGwG+xIE4qsJysYPJJLHaJLXpj29ljcnzz97+tsAtNUWIRzqUM1P5POjlyh3
MmsfLXAkOLoySP7Jj0gSQ6UIaZh1D0iE3CI9hpRqSCB2UF7o8bycyMJAEtJe98fqnfMsHU6PYd1c
Pvc1EzNaxfYArriFP/1ee1TIcQlR98hReaQsRGc2dWrptpzgYkDKxV4uRzIKycJBtTD2836mTegC
SzVy42SU+Sk8/wmIDZY9hUtdSn4Ac6kyNjV385zH2CsZibLIy87L/XplMlQH5FomBGPRzvTe7Il9
v2W+UYcpCCFU0fkYti03dCrkvRDKHOEL34tSpir0zcF/3ZDAQ5bttX7yMgVCtrBAg6kWalI9Tzde
NfeyHVLslQ3O+/+Qfxj48VQYUBjCpp4fG9EcHjc69AkgChm/FxztpO92Da3XIBGakMaazqxm5Mb5
6AI0l9hWjX+rjWFyEc9ERI8obFw2MS7d/fFjQmoa7TcCJ4tbF6wvE0fZ/Mu1X9+U2T30QBw4RvHG
2jXrBWAd9yHhhoCU9D540Veg+LAh2hO5+hkebfh1hZ0ZuNRwsktPLpyRRVzqhxFYq9Snk+WT5EPJ
wevtYdrnP+8XgjDox/PnKva06TrTwVtuHjsDPhTHT8xK3KMLxEeSK1ldYKLLuJQcZN65BMlmzx66
4KYBIbhNFpeytG1pTQnC9IjDkpjhU1XpNpm028giaF/XRwNsU5uAFHPfeA6QJGtJG9QNFKqVQhT6
adWqpqo+vuA482RpeDFv6t35DoOtiOOBUUoyj5Z0ERafsquBzZ4zfXSz4cA7JRdNqws1OAjsPEd4
iCms9/CG+ioKAwOhqwVOKQtMqCZEQtkyNG67XI4imQ70cMmBovWF9vJO9i03BGUtl6plKAFTiQr+
ruqZhQqsFM5A12UyXmLs6TwHwcuPH3Gc2JAuyjYioH6WT9GVrnOOVkAKbMs0ufcthtlqQX7Nd5ws
44z5ubkSMEGyBY0b40iG9KtP0b3m5740Dkux46OdkKddDJWs0atpdgAuAi9EjVPp6bpW8scIqlUu
ZDC/Hb3oC2P8keoxNz0dvPZZUVsFcYIBk8xXtv7faQG9AOc+eXpvFKIT1siHBIX85ghP2pKmtBtZ
Mbbx/VUA9HZ0fRJF1NZ3ehytMb6DRyWK5fPjC6sJxu9c6oqlhLL+9dcanUK+iIqiEzUAZIQnw6WE
maoMfb9CNZiUS+QA9mDkBsRDmW38s8Wbp/Iayd9Ug80mEh9qdfIyB/1LUK1xJ8HK24SG/hEIvHif
CjPds+rrf8MDVZZs+eiXRtoos103ep3TDYRJgjqizfSeM8L6e5eAhdbM21vxPzbGpp1K6bEBCYuh
uU1PwtN85LUuVNMZCnEVvufzJrNbKuXFlqDqod8jdW8aFpB1RopUU5fzM6T34GTQg+/cMWb+z2cm
stX0A/xVhw57+4b3j3GeY/K1LouKqruQeymZ95qocq7M6kxq0mrCSI3c4Edkpap0XIym5ISer205
GyFdhTaMD7/LaAcLlpwmEwhqjgHp8Y+QHojw5AA04okiubRbeydrYQrcnVoGlzMitr+rJbjPzcQg
A2YwBHH9qL3kFuRXAr7z4zQl/UWwF1Nwe0/z1JMKofkNavBTYQEJydhcBp/XQh+APK7Hocw3KYjt
nysy8Ipy19iIv3gDr5JieHK9LMp8KbpJXOAcUnAE4G6PuLthO4e+ss+pr4Tv/frfeu7DD01V54Lv
CKTZWzwuI+E/vDqnx2m00kTaYlDb8y3Iyg8Ryl4TfZO61tJDKuHxyDeosjAh84qoZWTmZJ3c/MjM
SUQ4Z21cA3JDbklzn3oFopUu742QKP5EWBnPce4MwMBN77btRVCnXkcLWHRlOAEgJgDwvmXPPRKl
JPbD0thrBx5AfXQdHrRHHCeRz/3yhZoOG7hwBjiz7DZYHN7LHig50oTm1/lZGyfHIVaT+MTnTpO7
Ei87ll9qfmyPq0T57COoHQ6iF7D/895HTjqKStFWL1FuRlgXCAnNHK7YrFkluVN6Dqx2d2535i+3
sQHPK4za77BkvL8P1sdIlSS7PpSlgU50zTejqcPSK99puyHnSc9YCKueYkDwuHc+dJB/7pCP8+HI
olzRT7CeZVDVqN6mLT5VMQP9d1rktfKUrpRwBbrKOCtntMdpSr0IR2Stk3jJ1zTcvfsSIKPJebs1
R6ATxLgd2vj61/au6fzQryLFZu3tzHb0dDoI8ul8xxvq0VU2fJMyuJ57ueiTVWN+c8IXk9gkAmza
w1WvNYLQKpqiqb1tS0m/BosjTDz4dY1CjRAmAfEV0Isbn2f19OgkqLpVWzLwyBkCWb4h6DUavOkG
8is1TRGLE3zwICDrgfiHlIJWPJVvjWdVbM6l24t4J5z2MTK0KtX56xwvuwTZIqv5KHD7+Y25vYLh
tbSY8tTckVpnxPpE9jz15Cs0DikWzOsCZYMD/Q8moTrMadhmFIKzzGTDMvtmnQJrCLYRiELr65cM
e03oPEvImwVUIMxIfvzqntjNBQnH7YBF0yt7gxMVVwGTMDTZ24/Zstrj76tCjKkROnPK+2nxOX7x
TwtPEis5UEg/4ulIb942vmNjUgHOWZuuipi3chOhAj3hSzwtvXPJOPcN9rn73KuT8U8WekN/Irai
+89K8Mv+NvwvEX29UZ2FdsdoBuFzaRx0bfavnGUll2VAXUu/e4VncM4g7j4LAcnTd6YYkDzMV3hJ
vSq5aHd+5+kHxo6O29Lkb59cwB+IMyIlLYVR7ZKbm6qT28HXNXAk0vMDhWFcRn3q8/cmvTZnpfGM
+HedawjaOar0UyjiS2PyzyQ6oJ7RxEpdGsZ7t2DmfsVqDRhXABmWtkHfIUC8uTnAdPiLxb6zY5H2
/8VBqMPz7dDL+G1S/G7qbjepZiWT2X7ThVw3gfWWrIOOh3BPY1GQ7kiJuvn0zofbYwn/Yq4iDptb
0rY5+coyG4qqQWYtWwfh2V03xjRwoIfOe+qfZLO8p75A91j3zAO3PLqiYfYUiuZ/KgVib4HkzH43
uK/UtMNx9jhGNNfVumnijW7oDvuUMlpYoyUfllSyNQsQv0fLEZCm1K2VW8IS/jm/WgmrD4OBtOKW
I+sxWa83QjQvbZfTWj1QJy1KfYwWqJHqx7V+vipRfHB1y+PqksqcHvb7v7fSyUwLmTPwz/skFhxQ
moTauU0YglJVkwcOgN4+5toor4geM/yX8QOXPbMo4GPJSTcyLVXg3HJA4hJ2Q1D7voiUIhPzI5fI
NZIrLib6hUwdlvvFl9POB/uzLjEyvGTKmXolmkkb/HGELVcGggZMs3WtnLYenQn3haZ/Guv04w9L
EMSl+Kj9wBcUf5El3UoK2LfRxXXNDcln8V7rJ0AXjKLWUzKxNmzYRHxbljRNp/9YOtEcBCm8zpx0
pnPQYZ+rkSkYaHLh3lbJWF8gxpbtRD4+xbNjH+SpPeO1E1DdanW0L7fqP0owYmNKU5rrqzl7n0RR
Xs3Cbfgc6A16fKmBze4oW0Q4FNfvwvrkR9GN+XYAIimQwGU7hH+ccbd7TPuMGAShaM/pSbEm9lDk
A+x9vqQhCjtjrjX7PKmer4edI1EJLhpAOyrRFag3MLsuMdSNOL0wbnoVOhQwj/Yd9KZtJeYzWKqS
e1Zf/Cd5fkKpIy66RP3YsOkO7Toi1nXHKIwBisxFm9q75g9158PIPIhzQ+zRBDbNTgravrTMAOEu
hgjvcf9zaY+Vb7Vdy9A2yOWJyO7QYIc6FZsxaWQPCjYFw9xnvn726+/VS6lxNuCwQhIzil/Bo9Yc
QynMKzvKtHL8Tt4nOsNyKoXp/zTP/jPiORDi2wmRiEjJT72fzL8SWPU9sc0ChTdPCa6W3MGDbawO
+X4n9JW3jp9kbNv2xo6WqBFMfv0Ly5LIOgjgwoY1S+wIlEKZLxNUwitMJszPFL1g43rBVKpPf+y6
PoPy8R/IGV0WqB4nQwHsxlW76RRXs31GW63kwHiMErWoSnLN1abwvt2zIe8xolIS1kYutXmh0ULV
16Kh5/J/Ok0ouVGWbzTiT7mCnFLjt6EXbqA1kisRuuaExT5QHvCxtW7bpGZ/Syu5k9U2ZkLHN0PY
oOKxqTaah90M2EBmY77bSENLUifZ4Qrf1t7C2kyfWMza2zSEFq8156N++KRyKkOryzS7eJOiH4E0
80l2sAy9JI+K0K/OKvQL1Kp1z/ez5itLvYQotjQ/CFsRv4FaRW1u1Lbo+ZLr4wj8+pQx0ICc3edC
wx6aaVbMORLM20suIu01o9b8C+LqLg8SRL1dHLg5/hlWusDsre5+3xBFKBgpSJgoWucH/85ItAbq
/5qFNbNyddETabdq/pU5ToR795zctf7qqVe01dopBQHQar2WUCu/KtfwJ6TtnGnyDgYmLpGuLM6S
9W+c/2p/zHHiCJmZbkR3zb4Wiou11iiQqVSqEfxjLaBA6uDt0rnDNLSYl0R/zDpQNg5QKtG4n+r8
a0OHXCWtXdwhzYqBmzqsR2cPJb655+7q2uqlyWgc9jyChKri58z9dAQh9/rGzXMVN9eeYyeM7Z5N
a6GCwc+g261lwRhssBJ3EGmB1G/zDXyd50feRylsVh+IM/XfdW41oveBULfCD5CTbNilVi5nDZO9
muUemGDdP287ZhwJuxo6ZeattHUmiKLoTUKChj486YfUDQqPzrQhiouVtzbIRAU/aXzu5MUaot9b
rEVOEz6qXawHb97+MKp3kXVwfn9LSNwM2dmn2ptLJl0tclsj574mScER8DVPnCUHL5tGXYDTRqzv
18/7w4dSuuVgSH21f4lplaIP4I3uq3ZyxtabYGZI3TfsxQ0OYd46sJpRrsaNjWWSSyz7Njv6pnGk
+6uYhp0yGSJnCLWRG2b6QHhPyXx/usK3Mh67ABmNqYu7tuMpD5/HeDc2kordpgO4yTg39IHdT8wB
iZYXW88uv9WA6Hv32wnD12zvSDU2HW7S3Vha1E2Bgxmxq4OksxtfatS87fXLM7EE0eC9yZpqo4f5
6/kG5pDK+5Hv1N0QP46RzKdFB0fNcrvtJtNXFNUMMrPWxTUsns/i1it5L9UE1Ap8leoEMxXbjvYP
0rG2LJKbWJsdBRZ+SGfQPJPe5sKg/6fnJ3ZpE8wmSvkeTGbtB/9mayQg1rnD3aHZohAc5QCWwR/b
ZN3ZJAH6BH5HIZeYvV0+UNNZA6QbzEX5RW7Ii16NMS3bnT1N0DUxnWnwryPh2jLSRKJ58MRjG9w5
okDLFgkigD98/3lCg/IN4LWJObnCdxCmm4EvDbbypN6fxVn6yHlBzYXaXdHRrbQBjl3ECY1G3u2w
h1NywWAw2Ucn/sq8+mpVfl34d92nnKJQUDLRcjso/9PM700HKYYBo3UmiuM3GP08DZ7GGOctjjBd
PYpo53i+VHlqTjBSTWJlCaFi4TJILWWQCZjjTuy7qylZMJ8QcGRops6zF0Ry0DWcydtFSDMlLMY0
/Re2yZ744249gnKhncjoZ16JcPcwDP1Q74/t3uk+LyRdVAS66Xggo1RLCyyURZBxbm//NSu1EbQF
t50Mo0czf606DKZoo0aot2P42CLaVLkUDE96txXFEqUy2iliqbpQ5lm8sS8IO6UsuT8Ruv2R9TLW
skSHmJ968ZIoBa+zTDo9A93bbgUjHn70wGXEWBoSvgAYeAunF1t2uNySCUySredPHyNx2TzMNK97
GnfGle5dy6/yC4GfiFylb5STygc3Be4i6LwVM4AkH83aXFMx+zxeWkrYLWmUzO+9Aq8OlRfxmgAQ
oubVpFRrsi/QhtNC8/echK8usyeCtuLeHay8gS+rtt1los7eaNFtEYNcf6qiT/HnxNBs1Jt21a8j
SIgyw56+1OaT7Q6wFrhzFz7hxLuNPFqmwhiqoxTs0tH5h9XDmjHQZ1/d+rOjQciWxw9tsDqS0o2c
JWLHUm7SJeMpxFO6GeNZF/bNPjibYRw4v6TXJfkwmyoPQsKCnVfrgTPBE91SAMKgHb/lL2G528QU
jCO6zK1pyQYnRiH+XXD8XeQYA38lCn/Phqwz8YiX7o4ZcNlQjlSmwpAkQ9O70vj7HLMVnkvgI30C
b5xJJDTeC2EgNHnvvmmPeOr1sOUIIXu20bVdhSTJ8dP59ArBEE5hNE0lLBvEllbbq9i8bWnZy28C
GxFZI6KOtR/fs/VLnSvWumwq0VoN9rR+7MGjRdK6T9YDDNUclDkrCp0JtsfkEEJWzSbgN5GBDP4P
Q7Mcct5dSq8vk/tRrVzK5J8U+HDHNKFI04anZegYdncfO4xC468zrxOlg8Ojd2fW4gm7djXccqLC
kmrDeDj+CuKXhzK+Z/RqAIDr9FzcLZdpVIR7tGihkC/QXjqvVoI/bunVIDRzOcNDfZfo1j0dboLX
O1I0JMchd9K9p4iRrshrfdLgncdpiW0ZmzuevxTtokLKm747vrP2ymJW8znDr1MMggWef2XY6QsZ
T/Iu88hJ4z7jn0vYchvgk7+2BP5FxE+uqh3v7NJbG3fRIy48W30DC3bN7V+6PaO2WM9dEF4OKfjC
/D+oTuvycZCv3zpvKSXuS2sibDaUO1cNddKCE+zVMbeBPdkyBdDu+GFrc5Fi7miYWxuXDSuswCAb
oVH0CAr5s1NqDxLiTYQCXd8TeUK8Yw9I65RLlBuQJIEfizqg/O9/d9bdoJq6BARIcDSaDIIw+LH5
k3tnKunhDh0RGBAlWtNHRZqKVs9RH/TZulcJwcqpCVwGktcnHtTOndisuFLZqZxz0tLKW8/yu6bO
f74Fa5fqvpRzb3GmMMOYgrG4xQQXCjMcPFakmklyCNaM2f2rI4rLN346ogfB//VuHNFncOmCEG+C
KmTdWeCF7wVjFU53BUDlpVPS/w/agjZyQ8eUrIvQ5Td2RdLsj2NnH1CmXRMHtt1CZ9l9CZeqTU+D
81OwTcBo3Ng19EOD39d9Zn3npswYcuo29ZxjNftIJPka/d3u2waL2HVAOttAQkRQqST15Yk2BuN0
O8Q0E+oNdLfEm4JIzn8s0Wj8NgxQATQb9jD/8zwXYFrf9Mhj+c88utGmG4108pUeapaV2Z866DT5
hnyn+NQrW22flreY5lODX+P1vCZQ2yczBSzt+gitX2CXSJS+VzHYZ7OijtLTkop2QdRfaBByS+FV
v0x3jx7b0TQfpoCRxiNIz9mhf48kqYTlot9+jrM2QB5J9+wdls1t0OBNxk1M6ZHXFRM/zBCdLotQ
F+8ZgnqLB8/ZKhLYp/2uUXHCu475TzmFru+sDJtT6QZKH1seBoTrHHzqIxy3U0QoRclhaYpy+xPF
owwC7HrVHV6ue1bOpYpJIdapYdGr63sQRQcrfu8fbQaORGhIqc968CAGMmkBoW+lTLtuNKN+G51l
jK8i74DryLhHVYAbYYxTLdOoozxspjCKLuSlLQmGl/xoxsNb3UcxWpuSugd16hu+06sAM45OWSKx
gBXw/CwVBzLU2VXs9nsx8oeF5f+Mu6eyl4/3eD9HpFLnkwDINRZOeNtD5Ef6hyC1dHwt7MGbvjL+
/qLIVN/IdwynApy2wDjXf79meDYCT4qbxHhE1aqMuBHCokZndZqqlj6GJT4Rydmsn8v4F9j3vH8p
O0RSuNzpm4rfaWv3hwkizSsRJzRE3Kt/wDJ9m45i6aZzztVTp2ndFKYbB77dnb1sDhuQho6RJwGV
SOCtbQwM/cj6bpmrpG2nyD3SGwG7UWllasUnrEJ2d5CKyHvCXolVh4RK1AGDXgtq4qP7sfcnkRVQ
3QgrNCC/bCxd+JLbUJZMvYruERYqM45qZsy+dfoBd11PXnPQSD51eJ2swtErH8J5EoReoCPj+KD3
85nVdc6O4VsxA3Sy/F3t8Vr2B3h54BGWC3AIUEDK6AbnyyKwnTaqZ/9uvT18BGuApEKl02u9Luur
+FciROGsOelUWISq5d7xWsYbpoAY02ql+oo6V66Vp2qH2V6raGDG8CI/DON97P3wdjYKLKXPlE9J
755rLC/OV0F+lpmqRiR1lX9rPHSsgv09Nal3iGdSRCC9dvsbbb9TFgMkwfp3CZQcxA2AyZbTmzuA
NO/rnLk6ztxeoewQJx4XgEw3p6dPl/vX4+zL0VpE+uM/LbbY/ACe2mYt823vB5HD3hsnWOwXW/K+
NGCxWxNrNhzCC87XJJmRNezU+IDxZVwkKbeteDDe049O9kUWucklrm7KulvHVsbAV1HtHfYC2WTC
n9EcWLmOamVJMPcFoB/kMQWBxehW9ffOWI/RTrN+WzwyPSNVSwcvC+edwo8RXaQbMVgoFXbpHym2
nlgRT0cHzAmW+FYW9G5nCN8vShY/HcNa+JNj6TXQENGpDbdL5FmHEZQz4eZOyIACvC3v0nrA0pPC
BIRhYh2jn/DjUONK5NSCORJaY2tnjcYa45aolzHllrAHJyX3B3gZvb3gV36E5YkdV/odlM6+/olL
ZjxT/dhaGzlKItvZJF69PjbUP54JxVnYkLGLrRE8qyFbF1yvQ8TTUViVSxDSVMqO7UGzd+kh5ewa
GyY6sFF85lZvK2aHP8Kgj1VtDaH1FWTqYuC5S4b7+pj4zZ+6MFndxIauM5/YSSfOlZKRJJnW+Fdx
tXxsnfdPpY5zijG5uf6qY8+vMn/M1GwWxgsgyb7V2zW8AeKli6PUcsmEu2e1+qJFqbQI/P84faYp
7okhY3UFaTxj+mku7+3LtVTC9QFx+7RNslNTUAu+udx6pP60yz6S/px+sL0SoPNvrdZWfYHKYsx3
jK+dWWzD5C/kNJGV1VeloXOL5099SIfSh8sL6wdahpCWVV+k9daAhB9VU7Is8Qpa+xs5DHPz5C+U
ZfE+dIOV/KH5bFKm1GqbMOUz0/STwaUVnBLGOCi5RUk+9an4ID0CdCVJDEESi459vaFxk4ejNjTn
IM/7rrfc/oB2Q84VUUnkqmdEsSkhzY5B/CjxeDG+pd5/uFp76N+eu54LCbJmRHtRDwauKS/rwuqc
0SEQKSMxFIfqY0VxgZSmPd7s/abpWcmH/3tWVDs0SELvQJiVeBVu92rVXQDxzqWGKrq1fep2ocXh
PUCPYxIBSGtD8gyN3LynAvBvtD25QPS544VkkiFpzLGsRFnyrPvWQGTYzj7vttQBARAdd8ISRYVK
gAtT+69IAwv4toz//hMkP0NZ5ZmsXGZ3i/oAQQ4yVLIl8u8O7cfg1irwckVjg/VA6lu+wtDmIXgD
4jf4kJAxWe64Rah51S5Nr7tt8/zsH82YW0gnonlVv2e6yu3NVB5RsnvquQOY5k3l7TAPSSjV2kgK
CdPpodPZdhTfSctYsxVAX+ux7qPn5Bme00g+qXs7SbVwV2/jT8VPrCeGyKfyTZUdqJqsk6gjNUCd
8WKwfYu/O58FVWMWAPDg7StCwTHmmyxB3How5AFbEH9nDhQW4glj0mz9xEhCr+6sn+YOOlXpLUeq
jBM8uxmc/Or44cqR/sH+hNrs8s7SYf2FbLON5VKzo1HjdtgfMG1D+eGSWuXvd7p7PvorrO0Fx+Fq
DWygJHqOGzWckLdV3m9VMhEJMnE8WLGLtt3PwJKoqXeclDGULVnqz+MVA1iwDwNz5M2k0IOxtj/A
IoUOO0huiuaTRfXlHwyya/uCd1Y4KnUyKOHSjnWWDB+31+YE2N+67qw2RVnZzhK7mqowtik89lgg
FD7NZLh7dL6n+i6N+KaXyxrWpVbKRujFQM86cdy5mkrDMHRA9zUKdbS5j1abanMx+ZHo1CWBld6q
vOsih0ixrIwNG3U2bfdh0cCb/5ETQG0pKAjE1S8s4RRqJBUKyjsOMjKTyxDNRtoGqtjDX7WNKJeT
hKL4AAwrS89s2mcC0Vx5z8+HOdikzL0XTK/JRDovYiRqJ/7ssJ2DOYxC64EXNyRP4BbuZf1KS8r/
SjdfH1VfSFOPkqZjf8Sb6Y2miWXEtj1umW78Y2z211PXpdQtODiVzbt04ELVPmmCBcW3Rs4SU8pt
1+fkKBhZBW1AlD465w4bTsSktWIhf2Vy1lCFwkZaLVQ0ud4v8W5vWdJNs74+Fvq5DTl3PCyTdoGc
TbaKm/ggeJliPIXEfKz+8zEr2oLvnB4YINQBukCJAs6oGQsdP4mF2u8v8JVGz+1VL5piZMbOwx17
5CkIkyCNBnoTwO/t6LQW1k/DujXIdKiFZIMBW6rdNzu0WOvu76TNW3zcCHmtFbvAjX37C1YZFCnr
e2KAsbckvCvlPZYm6JhkzTUJynEs4yMKYhejSyfax+CQJGwvagnlxQyIOueP9NmbwySoyDsFQcH5
xQjG/lx4VILGRUMpVR/yca7nzDP+0v6b4btyVDWM91eIdc5EoftXTWErd3wx9RC5aI3OBSW3ECfT
kz/FsiF2GKG7L44YJBN0Qopzwe43w1Ol6Rh++F6OjrQi0owB24Z3JZ1BewT7z4p8gtE6QMQdYFAC
Xmbhq9n3crouTZ3wcZ+GgtiH0VA1/pNqIL3YC3R+FOh5wVESerZKyB6VnQna+cWKld3ImiiukJzQ
ShTdo9idUIozis0U48Otbx0xSA48HCttNy3BruEyI7izN4UbkMfRggu9oHvN/8dNZXNjCPFeHnzO
pz4DKWarGtdpy56bKGaDtvG7wohiGCdwuV3SDkhx+QxZsFhacAre7WcbXOffAdB3Z4cr50tJs2h9
QlvF8Ihf/fTlG0P4t1YqELb4iXmtRW0yhmUE6NPgq11WfDaPoV3JDzDyrVSRqiTKiSgTOQ3jEsF/
9UfxL9kUXYv4XNZK8ffqA5ti0sUr0WQqAQAA2RL7WmWt826hxlP4nGBZ+7bK0c7x/3HxIN1X+nO1
So4P1iZqmPYjOPnbJbyVWNP1J1b/oDjzmVQP79U6jlOZ8kmQsTHiobtWF5NtMlFLKMfu19Ikc6dJ
/J4R4cO+px8GBP+lKOrx8qyqx6UkJqSFtfGnMLzGBtHD6iYX2CLyvux/QX9u5+U8jMM/O2diTPaN
qIH5dpzhIyDZS//WyJIjhaBju7PPzEzmgfeNvk2jwxACwkEr9mInyrj2VZK8TJIlhew8Mrzrc2qy
MYcknNtcToPzmQQi/I4l64FythwDmD4f/HZPv1w+IMFqi4XIeGkrFElTbalyk391pay5clXx6+gw
K5ic/R3OulJetZTL64bnRwR/GDP2DF3Y8Kf7BHx17S3mXbP4KC3stHkXiIo9PtTkU4pxsns9kGIS
G1oh5mw8OBQUtuqemv0FbQhxWwcukD9pLhyLJKRjiF5I++gXWlmtDM4/68mBrua8g4D0kAGQB3wk
M0mkcGQ6EkXN1nrKO8lFOiZkfHPkGMt9ep67dlcsivsEY3tzziyWgn5pZCoDBv9nebhSM/5vjdTG
HKy57LDVxXb7XV8tPAUBwXWxawhAqW5eYZWq61y6hL/wtU/qpvN/ASWA5NEO1OFfnNw6ZHgak5b/
EuSawbhzWTeWJLKGGX7efl2aM+0WNxG04Lr6qd1qyO3Sx5PiktyqAzhxZWZDEOjYNY1+oWQlKy5z
KVXrBZxw0j+vL32t6uyI2aTMha8tAT8YR+d5e1C3wug226x/irsmCtzOW+sfMGWo0ba9ACWv1X/8
lqIwboXvVqzEN7eLw5dt7plRpcYfnF9xA2HlNfei8FMy0Yyac8HXfmaul1z2s0N2cXI+R4s4hV0G
SIdOQ3uyQBdLwg4CVdozIFZ8W8XVBjMA3R+sltdbuOsA7xu+XleDm5W9QJadWT0z7kbezOlf5TQD
KHN1gdWigb9ptN+uyX1MYT6AAn8/GI/s0FUf4+6+SuSvmef7992SmVD5Wabo4O36edH44TAzji0+
Dm6TFSg339gLup3KHz8ay3BvvsysHRfZq+Qc8rXuWl6JU6WyHyE2YxEizWyLJgflKaOuLCOg/BTw
9XdX3CgnWr5Hy11179P54m++on5J8T/Ap9XnFTdFE8aqQme5fWF1qZz7igtFsHb3vLx0wPioiZ1a
J9devqfpdhbDy1CZspZ+fEtO3zaSPMwp7NLnkcL6MAYBtHTVJZDUQ+hTC3xF1MThFNp6MlKLrrRu
hEm6OHrjGtOhGdK0WpYs7BGh641d2yjeoHKTJXMEWNohFnUaZzCgQiD7tbFYBRU5YLQ57MB0k16L
AM9R561T3QCYRkBKq9xBjc2mtm3mNJgrIehYow9GLkmPlNjvuOwT+O6FpQz37UBfWf9Mr9Qgfus6
tNAJP6NPKsJZkaAY9dnBnE8Z7MknF1qq8vr+GtoXGRv10OsD4gT3OtMOhU84hJaHf1PfXRb+yp6l
So+x3JsQI/lfzebTCd8QbJHetI9xBVbc/2ijW1I/9XTNYZmTZ2kdKFhxHLJvYHpRtvlQtSoT3WOi
IEEh+bN9ajhMmMxtc1uqOaQT/lrj3HgjDDvGj3AWNEw/012QzYbBdxyNEDjJHmzMX+fTnTg2JcWB
2R+AJvyv8CTFAh/qTn+yl3DiEmaaj3uaqe3sn9vl/8TbHNqrWLg8z6jwSufS018Dky76pimXcPMd
9Q9L4H/X+Pop4K8oY4sM+p6jVNaRxH5qdaABcdfzlBmLOp77puXLVDpUFTpEgEg3VJKUXdt2sbuN
VMEjwtTsrnZhhUP6o3VoK4oxF1bljucak3qpqEodp9b1Yf1W/jvK7o4X0yP4cweS3Y4YyT2kqali
18j+n27p9xuBMFIGPorY9ckxi/lfRRfaAQdVn177nGA1OsMA1UHXSS/bNjG26teeLlu425xhmaRJ
RRI5Zf4OyAPPvGWVyFe/QBsFq0TLnoo8gYacyqidhzRUchpIVkYxs/KZe5CdTuHrCAnzOnMWskgy
m0FYZVjkTEEY6M4pUuctxuS506r4J89AOE2pTOhcJLMZgvtoYrJ2atE3SSMQGR2/lGMnewQBIyNY
VO//wS3LLsFxlSmpLYXft1Q87gJOFM2fG5gt44NnkYpkWD2lqqNL3So9a9M5CRSUUknCdIn2tBVb
EL+B3vtD8QTzZNwLD950GJOotay+87TOKQ9pgxkT8AiD1U7SPwhwtAYTnZurkveq1G/YZH7QtZOI
AvfLuWKwMILn3Fzmmy1G9L2G6Eeq0ZefWsKCMitJ3zh/vx3I0XBxB9xV0L7KGZRu04VMaS/S9X+4
OsjH6vo0FN6lo1HAEJwB3ZQU2xfyaN90Xn3ltDN7MbQeVDT44rVjrFVWYTOzkiLY3YZMZyl1fPkK
gRK5fQ4IbFk1mF16jLOZIpomlkwVdfmOd4CvGt7B9iPjwWhpk/7vRjMDHZeb6eNm3z9Csznv1HU5
jUgllMkpV9y2aPWTXCco+UlcLgoBJ1el3FlvkJZHc0XXElMta/U4HgoYsd8e489tCLTW3G/CX9co
I24FbMZZ7WnuSY746wj4RONvwhYpSzZkm8QIfBhVUiiDmr2JCzS8FQ2PUuMGgQ8EDktgy7GplD4f
ksUkHnDDzLjm+LmiXQfahQIIbU/C00yUoSqjdAVHctnhMjymtt+Ng5z4GIOcd3xOhj46nufAhLd+
LET0MPIj34IPHd+9XhjTGxJ+k2Wz3Exyh08X67TyJCalByenAq8RrpTtJUysdb2cw3BCEPS6REJv
cHJXfgBLVsPmiH6Pki6YCkUliQxjvHJub1C2io99283v6BVQsJsmiCg307kkdTKulUNlfWdIO+jv
hd9EQcnuef5KruQfGOlYrY+cU6UGQesEZPreWWYDm6NiEIHZlEzrjXwnWMbp5hCZ60CLVznUxQty
fl9uQey5U18aNLXvv+cgTCi4dO1GDf0HsEF4Yo/+Xo2jIn9B3qU5fVDOHQkZ4ZxVTY6nOc0RwpcI
UOd9gXSKg4xoWaqfPVP2hsbPtlvJtPLk1bRo70Z3EPKgItqkm9FjkOKs3L8CPaPP1DZxAtEyZxOt
UMaH3+XSecf3/eIuwsAg73cwPbGvV8EfJP4BbMvLCzGfmIx0cJGhYDjuBnuzfXUApFuxgl1Hy/y0
j9kP7bpXwXSLtHs+nBRpLx2zLdRIWfxHBji4W2b05NdP2iLQVslm8wdOvXECVgIi3vRy7Zdqz2r4
1vX13DhkbuLOJIjoKGsN13Od29k16Fn9YX98XTV8OXQ6bLLUQmdXDFoaB8ykxRdPmH3SCRJ38FQt
uybzkwktxyw3kzKS1S4Ur6fmkYo8ri4+IZECcflHptYLREntgRU7oS6cwjeIWYje6XOl7a7F4kGX
RVgBO7l+V57zE2wS29sqx5Oee6zoy2JnHwHg5Im9NWKrw+N6bhoXGXIPEn77MgyMuRBGKuQZHWEB
zFtQxHGyOej9nj8m4Ec6eLdDPiVo2t/rge4g6KrxGn21I0IcS3wd/jE8OitG5nm1e8PSJqjeZo5j
N51Rd2k3uDqZeuhkk+7d85B2vJlNWPXL1QYPH2cnww/KB4BQSX6CnZ2xuOVQe4jgd+DK32SCjPwa
a/WH412R7HRYdTcBQSUHVn1AinxNNFFmEQnA8ljrTr9v/tPPfNRJlC4XcPjG2qCyOeNZKU4jNy43
d5kGXvG2d7TcTLwnz1foL+BDbZ3aB8XQDhF5mu9wVcbQa/vdxtILRmzWzNPXT21I3TQFp7ZG1SNC
kX+s8BYUrNK9OR0yPpbXLW1qY9vSdFzO9c4xJB7q3QEA5YVFiyicm7iwOOYRvlmVSjEvWyJzFizT
HfK24g2gmMnd4XHyId9yzgbAldKQIY0ud9siiZP8IaZebtvB4wN+c1MAetb3d94MrZoZQJ7JfSTm
s1+/7tiJcoG4NJgFX7UXbQZWap8HIM7xZeQ6HlLwO5Bxpg7slUA1Kp7uqZX88oHagxPgO3Jgt3ZF
JPWz6qsvoVjhexBZK81ksFeVWJy+Okpdz1VpF3aB4IjFs3fQw1tI8+7hiXEdfYqxbOwI+wTMOQ3t
ojmPOL8OrJKdetwSDifFPXFF2eN9yJeXXYwLu+YA84wWm0pWlczzxBX7A6mcTBlu4DD+04ovXhQw
7TJOsm1Nx69MqRmXCtqAdwGIUFZ7nGtiWxxIviVtosytRjmzz+qhgPI26dsVMaEp1YXo5kvnik2b
wJRK+w1A3B+iYVzOeJ7WmLv2KQ2z5ODye9IVxDR0ORdjgKH/DosUd8yiBfTRMUj3BGa2K5YmEnWi
VVQ2scIAwWyMlQJWwGGhbHulLMRGzu4/lZRxc2khxJJsKNj8nIhk8gWwyTaCmuU9+5Xtsdw1HZr4
tVWJWrOzB0tWz22LRFoJVQn6nmekeLMs8pRCMMxnrFuSVU4s4iFvp1dWMgBGK2qQycS6HToi1eJk
q0alvqESdTqzcVLcnh3LYxeJ6IwHcMT1yyGMqZGvDvnTa4xIsg4DdlpbopNSypJcM3effttw9WjA
+ndOAP2C/oRImd3y5YK+bAYJrn5daZwg3Vd6SDJEuPNw1KAOQX89+dbknWUFbuLhXPVycPjc+bb5
ilvKrZrXlaYD18/cfa4hVuBWRHTitV33nReaQH1bfwwSo1mrZLURxe0xruJnBySSsJqZp7GGWjgn
i0+GWM+HYcwFTjkKDqNptomSfJWPPBIiA36Qx17x7BbG1VUBEKVrUfT6NbgikJ2ZuAsoopB1Imgx
4P7aP+uhx/haJkrTWEbgo3RQ3p+X+pAtebWivmEM071Dk0P9ICxA02Y9AoMRnK6HWbZz50WshsL/
RBuxeafnVQm93ibDVJ2wIA0HcAhQ1WVF1WBeLPw+wTAuZKujnWHqbsaa16ztFhiQMG+KPg65+pJt
4GWA0DTuh8Je7Q2ZJwnJe7BkcD0yiTQrKX3J+Tj8SGzTmLs/5XOM67SmI9IkJDrrXdwotinKmf9V
VHitehywxp8K837+HpR1IoJeJqD32zjieZwsQbP5q3mprGC/EeoFfu6Z8JG2ZcJn/AyZ7IA6Pi8T
MvxL+M9ahMZQbYp+idfG8hvBfN0yXprIKpxyWFpCmrXiuXLB7pbFcS0ww6bkzE5pCuFOrimbd8x9
2QX7YD0rpvIr38+Wf+U9VMkFblYUTD25EC1fi2nCnfNIF3cysi7mzLVwJYZY6fhtR/X8iux+7KGz
uu16wH6CoYAOzBqAx++hm1hwkr04kivT/Poiz9zpn16Vl7Vv5lyDAAcsuWDn9lkl/gK9RgmYY+dj
rDqdMj/two9yoeK+ImZXi6VKi9J9i3rXuyMvGIIEz7LCiv/KtFlj+iLTAB6o9VcbBrVqLUI5966z
X9F+CNlrff1WWz0ZLeySOTjYWg5Btqt/YidwpWyuuiivFJOy8lpm74DJwRYjuo+8yy2sAJyj2H2l
iFUCeVX7Ga4rLol8Zzpstv4DQUrB/Wlrx5ASQLBt1XjH4HmzR/I4uhyqFjuyJEp9hs+jra0zh7jg
vHFxNunRlYLe3ykofdVACqNTlsj3eeL+4PIMuFicgvRRlrM8rChPkTChZs7w4aLO43QzHQy43YIf
umGTuaMG6zGjHPIvxgdWXxdHv92OtvEVzvpuD2vr8RY1VgXkY62MrxMR6rkh0A67/OJ2DOJEd7nS
JQ/yAIwtT4QYngZCLkvo6JUAe/Ugfh/ejN/4QSCfDquLu/vJpHe+mjG6IBmDFqXlzxEfpWzVJyoL
+lifNB41Zyx+y5fDhmIOyg+XipzqMd902JqpeoxMlbtcAYd5ur8YOBDzY6lD3UEtnPlpu8Dqmp5e
vBOYEQ9JXzx99PPFbx3ETNLtAEgoawwnwVTJk+iXhbZnkcyMEZ/OJTFJ2b+Yad724dYRcfHd5/ct
4Ra+45sjzKcWzAytMvf/6Rj1yyqTCPnHQ1XhQCfDZoh/Z5qaYPjI31iYSAlLa7v42PuR14prME83
36Oi64dn5UrsR13bdriVsV8oT6GCt1LmeEBpb4SCX3uROx5K0frdtXBnIxEkPmtrtCsA5oZDHYVW
5KDGOPonovcuV1pgHi3PIRula5bn6XdL+qFN78ONy0TwrWU4LElTEGpRBulLZWBp2aGYfsYqaf7l
uE0tJpxoorJSAGvy8WUmwNnP7mpIqZN8lAV3owkbz2nqzvSP8lXJLBI/ZDi+/vlhIm3pof6k24TW
VdkquKLeDROjSKwC5yKZIW5B3C8TChVUTZajMIInS2f7SPXaWKEEI0D/jWdOnytj2aYF62eYS576
E1jo7O50xfHghkdNFMiOipvEUj5XCMow/MJyvTBXTnx8HZJ6CYteDX2SpKccbopiEMWB9aiHNyRq
MplkzI6+eMqqEw3so5cuvjkbebfybv4ZuUsTIQNRHk8q43R0IkSXWi+VcdrqGc640gyrY/S2d4+8
t1O0iy9lFmIS4kyunG6DvCo4SnNvPXT2BBkpIxT6btlbyZzFD8RJC8SFcLTNekOT1fYkT6e20Pro
1yiw+mM0Gd63W36vJrWc1322/0cwGcZq3b6qE6OryOmYctugb9pkDGp8qDbl9TY+qcx6Mo4X6hLn
XQOqCwNttqMxsJn4dhz96sg5mM2S87UIIDCaRaHIxp/uxfCRxQzZ4ij9ymBriFzuYQM4sVWNo5XY
ZR0StPkYdbQ2A84IDIi2OVqDSgOzCgWRze/eS60emnkiNP/mu21HOVZAyLyfwRCt4yjdW8N/+/5m
UHROcbuMPzvL7m4YCOSdebITPdaNfoapMmXwiCWowldbHcLTd/O4FvoQ9mzr4PV0fAejYdzSULkA
uGABs96ex+Rty8Y4Hmo0RDd5JiqRvDMe3xSWSxEjy5JpGU9Uca3Zsd0FaqRBMmX6kD9B0gBhEbdg
2FZAzS4WSwziVxJYKplBZa/B9YdKwwnN87iTS113BBd6pOsC2bojV/Fs0g0KW5ta26YRHJcRswxs
kfmrGLMXh3CoHmdm3R+dk4kDlA1/HPgfTlheMyA/uDtgnfg6iEp0NNBTMjBa+oKeguZszIUE7QGZ
pt9GMEbFTVpqPQcv8V4B3H1qFAkXCoZwVE8WSk4z/jlHC6esRDDFREGNL8HMn36q3iOzW0VBwT4E
HpPq8GjIJSCD/u+mNSPt+fYfrNDX5VI0vTQv9JKJXr0cOlj6IYO8tW5XJOIk8uoGzsCmX4hRWs7D
sfUjIBcyl0WVO5Y0eQplFGver2miJDckLNQnLLVMu8NuC0BCqiwEX0UvN6NyESdbcmMLPrE/bSSA
BUYlD4+a+g6c8d0MKRK6ft3fL5ttOJQl8pCaHTGlUKXn3zMU/6mw3vFMRGodPMmSUh+/8WjhyPmX
lYbM0KgvFqSkt6lrAh5CaUDdphwC8w8mWn+mfj7TE6RdYqoQkV0eR4m8dz0sHd0XTgVzb7GhCzUH
ONSPR+pqSk5wS8CdHhoCl6V2+cWI6w38M2/FvvoEPFGGmaLqteIFJHvyahf834W4JdLI+NgfHt/m
QIfQ/FR5t7csi7p732WXRZuM0dyHzNO9sPu8ebuFlimvMaSd1kxd95U9IcTRcqnXFDe8pOWktlkY
0jYpgEIGX8rrs5Fuuxqw2uf5UkMfkXW1OFdCEX2oitqpu32rX5PJy0zLXu+ts4db1s/hpMyjRto9
oAtiBbiit//2gA2BjgaCI7wdg1f/qEbEwbjjfDAcoqPHGWWVWBXQi/mHV5RyAZDdxcn7yGo5eCI0
c47+XItORh7veRxt0Em/e/xT7r57W888R2SiE+6kGNzC3YbJTfww60UrSyTB/68x2l9ZUEE9xB+j
g2zFw1iYe16NnlYklkVTe9SqeTcPXvbJM9bFXs4nrt2nF5iBiMOmB3CWgayJOzyymAwb/Q/ZyPbn
2WnOEXUSIa2r72j1GtYeDZtYAaoY+hbeb2a0RAqYxqZMliWCfgePg5BxnGRNYKuLiSUp/D4GVFck
ld3LfNs8eR19T41Yj9Pk+/ynkuZOAInR0Kym4xqyshfnY4lcKP9KQdt6bq7yYFLnbzarBTOllorq
qe9AOd7fkH94LdjCOk78RKyIt2Rjm2NP145/kSX+H5XCGCwttlWDCbT68Lh2nIImmtQBl72NgEew
hlCOgdGB2rDT/sSRTJlmDkt5KOiksMxcncDlrramiPljBXkkm3MK9F9PwuVm/2NP9v6MqFDNwOdW
HM6K1eDVs3c74ezC2/GGZeZ0X7GqhKKJc7ZVJucW8k9O0RelCsgbaRTjjg/DmPDmcj6zrXKlTWLW
H/1wAgWOeAr5sX4SGi80y/cw0nZ4KOgjOTYMB+BNHMa4kBVfKMTLwhj5nDyeETMnK5RNhKTrqka7
lsH9RdaprgerDOnTnIEhAaEFH4FRCtFuS7bgILZx5Qjv3JuE0JTKafxQ0DHO9uLoeURtPoXM4Azb
MkCqW3j21XwoUeyWwIpnrIyIEVV8Qv4PJtDrEscwactmT/MIc2jA77e8MAkS9YJJftWaah7F6bm7
BkGYOyyqwJr9zROW9zz5s2M8Wjv7UUyZsv4MngVJbDz1vNXBujgNX89uEBu+LR0Ur4mVeusEeoV4
HrgtU9I+Sk3odmtmPi5IQt0d7rbLHwf6ZekqG+BrYTpAkb1sU2nRZvNHlTC66rtHSgU6RFW9iO0V
40NQP+h6nsILR3rP7Zj0pBxLhCxXKya7F02ndlsJmYuhMGeDaVUrk+tWuw+NvJEXOfms6KXzOEnf
NvNoRCiXq0eeT3Htse8BMuOzVnp967PZ702IfYE/ZWuuw4WWoD8NMdSDSu5F+028tT19Ty2F6R6p
5j0DPhH3+FnmgwLv7siHPeoYFLoS62uctlpJ6OMQZIr2G2l2c3FfnNtW9nfK2iImth9XFRvASnO4
XvBPlz5FZpUELHS5mZt6v1+4QccFM5LDXI+QSNCetEaGSj9hCs14Tuh3D8oKKDTCVvMfhhc1PIjg
dFbTgL5tiDR8ka/zZa4DgEzr1PkAGqHs+QUyZKO3/vyMV1blzqgAVR1N9KebDbYqMacHREo6GPUv
zceic++Yg1yr9GlZTXZX4nAtudU3TFVkKK0R2jVjEopx4smcr4nMswUglqdO6eLnDgNtKB6/zpCX
+JsA2edMpN4sDDGRlnDz4bXVZdtMvL6RxS/y0W8DYJ3PMKEB7XkAcphlXXDwdwjbRBSwIKFG/P4g
v9AQc30LZJJApOrvQulTEBYltEqNplADm7JkrBav99nGBCk7O83gD4QtEqb2Cu9akJdSCF7oCoHd
TA+R/XM5V32Y/7ODzID9ar7rgTvWGQEBq1sSIp0u3yCeM5Cv7XCzhjwvURU8ndhEvR34OYg4KJk7
u4Z92WqTaB6v0DW78zcIa88Q/E4baZbbaKTdjuHOmKQP1QEb3RkBcjLO5b1MmTEjCh6Bc1XLChQU
nF2JRfEXD9rotejdTpYyDwHsqhoS9m2j+BOkzJiIziGLHYtmTIX1g4n3a1AEnRMreF36QQSj48Q6
Ys10GOIIQ2TPxuZqJ8ieNZHtXz1+YIz4E4aS9VCXMSPwI1iN/in9MuXu/6Tp9dxbXB7QY94yCucR
YEkDSn/OKESMX+4PCE10ye1dq39pJ2QvSSYhFhpRgJpdqlUvh1rmTZMlOs92v6DbedAv3X73E6j9
g4EPnzX2PJD/SCi7wcWOq2RYxZGg5uyqkhFNM4XbDQsde8hcOFDRwHI44XHM7K9s2Qt1CE602JfZ
ZxFYx9rlRO9zJpDdgB7E7jE3zRLL+FVLEw/qOdcXnNsZYD1EmtUPM+sTa15iNmiuazarVT4hoSu1
WfF0YFdcSnTeeGm5GCtJw4fVzQU/Owg3URi+N6xW+BQ+uVH88eVCewmixZFG2Kgze/E8aaGXB65w
TSS0RJKUnfUTXb0fIFKo+qZDM/g1D+QUOa53PvcB91AlidlZWN2qbN+ygby+8DTjPoFvHHdChTrH
SFEfjgngkqEGPyjK6elXC6BFovhUxJdb3z8UftWFtR+p4d5JyfSdCQEnhMw9RiXUewK/AUyo/Hvv
kVVslT9lnsjzqAhYjr9yXGJK/m96DeQWqnF7p1iPJvruoi4zB6cPvS9zavdQ9V0OwEwajK7fxpi7
rxjCUSiL9vm8STYUaD4JLJAvGCRTFIwPpRK1kTL9sMrWLr45J9CKlf6pJ5BI6perRsHWtUIliDyf
m9TGwb1efN0wYEchjtH8VtDaPj4TZu6ERDMBULA9mq+zsgAi1RMqYoRl8Oyc28D/oJC11mJeZ+Xl
v6eYEGOwZC+8OWw9k4NVL7MUImgYYRyC1ei5YP9xaCON5uK91Moqpj7GCTd+1+ZXaskOQFSmn4qR
jtS/qcqfC6NJuTTTs4YXts6H4FDIM7IYzK039hmHYotmh/HN2SvIY5nVgqxxC45TJu1qp4m5S+dw
oAl7pIe7swcKgSMw2YmQ3vsMeP9RkO4PYeI8+hXreTNV9mZfhuDUxo8PIaDe9umNJq28dZbgUSHS
CdLAw2ZqDtYeaHRYrrB0vVJYoBVpTEMJgmkEJfDY99uSi7LPEJSEOlhwpcPnScc9Nd8G0OWM7Ek9
9aSLrQunPEhR6xVqvwPdLhCAwT1KEpGZvGm8mRLk9mCJWTO5PDWxCVKvgxrQ1zdmi3/L9YPNUugs
0a109o1XEk+CNOv1JY5BWw4geBS57i1IR0Hh7APIHAfvlafgqyrU0+EefqGE27/gm9NGTrt0iIRi
4XeWFl53yAILqqWONMkrKLYxD0c83WkHpDmtnGVyyzSeIwydn5S9mp3LayWBFo6iJyP+ER2YXd8O
QxvC0NdcMg9E+9RC7NRXQxE7f2oLvCeU5tD/CL6i32Y9dzNHTZjfGloZVt5qJmcLJH5Gl/GoUGAc
2F/cJEjNh7qUuhx2cEfT4tM9eA4QNCAaMJpjSPC3RJz6mpVRP1E1jMazpjOzkofOgeguny4ucS42
PzstiDQq4yoYvqk3vbL9IZAX1SzjEVtec3M0aIvjQ2zBxVLX0mKUfn0e0C8egvhj8lRavX5Hc6ab
pymuKpsg0zTGKhb46cXUv9ZWV6P+BJK2VWfYpBwkHxKIS9jRR3uxkcxO8eOT6JyAuFJ/NEwFAS/Q
eP+ytaOQlL8eskPGnKi5s9zLNrTd2MOvKSl0hUnsfUiXkrtYf0XFfznqFVCHdIZSajLI+8/6/fqv
5Y6bkMUqK+gcOve4xHckcYkv6MmzEjU7DmQuxq9N1jL6qse0SFgud+sSDNMBgK1HBQksuRoAGK44
wzC9t8qCipGAi0Quv1hoHd8ekUM09KYjcUjRVk2Lsa0gTYtPFpBA5G6o/Mqz9/fvDwYiEmHUX0Ag
Y7fI/Tq1ZmFGh9lhtvi59e5sedMOfWVaYBCYDcqZHEfcUjPCc2ecF8eD8AQS/HE+ZoXKyFDNj4e2
7rIzrwO1Ks2vQQG8d5FW/R+w6yZzEOyT4VnTX4Bz7+fe+z0yp7xqqiPXM9kd8yKYeREo7JHGnBp6
OXAvX3TvnWyi4HNdckS0KKoK0pPb0XXziX88bvUCGO7rjsneesZhKHRwz72zC7td4SIpo91CPtBK
gxv6PEV+8PO7y/rjfZPDPGITEatIHzhPT8GYJupeZkYXjvbrO9F7usgf5wozykr1o+GTNOFdGttb
ojEpwRiO5utLE4nlXublWpeBr+uztyp4zUlVNI0QSWaxMKHde8Rf333gWIaXsu787x8DfnUxJ/yt
0dLoYTGovlfFIB8tjEPovVKptEXA0du0y6OBavl5G4KTMqB9qN/PdPKwbfnN8uvs9Td9oyJbe0qZ
p7O5qPULOOVpRt4pQO5DdkUnEIv9N9XKg5IYtSQT9Wh6jWgi4O6BxV93zfJiz/fe5NuiS+Y0xWhl
SOC4bcBv/38yl/XB9pH4FIxQYqlfZITCc5gl/dCihDM9L6Za5Q2nwWEcrtMnd6Zolgiwo/i5IEKU
OVeEH0+lMwhzmSDp4X2LaM2gxp9sQIgU/jSI9OhfzJFa7/nA1G4omQ2F7YuuhRcyBgIa6tSe32YQ
iKtuhP7+aNGyMBclL/XnDMDKh8gjIYvtWPB0pueyoBWYWAvwOun3P+sKn+CJqNEtioEdDcFHDx9W
f8z00IdTo153HB1Y8KUhwcGp1V2W5FFhFWwte66wmSkD2QMZ8cZ7MDVgNs83+DpAaQhfbqVhOxLa
FBKoc2B1UMPYfve2Q2Ug4r4t/O1PlY6wOiW73Y6C6R2ddMcslDQsjyNPLo2H9pNtto+UZjlcm/pn
RkFdN2ILdF0tHv3XxIVkkVxKkVp6Tigzn45V2GkloAqryHSIoBgYitFsjGISHRzAXNNzClWfRaG2
vppnOpsY2wyNTmTQbs6jQZKLMmZT82RR4nJh6kRgpMmQz0S3g3XjYReeGEnHBDQMxSmVUEjClUyw
tBouRAAQnIz1apss+f0hWaSsEbtoUPQYPojVrPFn6ydHEZ7QvRwQ2YZ/CaIClYIpBpRFkR7XBLwg
BeFDHPJoEUEAcJSK7yTqysnrryouqWclvKJfnnhJAyucO90e+tu6DvBx+1FEO1qhsJrft01m2q4t
6rGOCyySr7pGbg+UuKpNPPG7pTpSGKkVPlQe0T13zosxE6+uG9oxlUYt+LrdxTWmv25uwBjFOu8C
1P+lHB7LgNg5nmq5eUnYogXLKzN6u7V5UzMLyR2dBXJ6UTsm+TTWkL3qA6S7F315RayNpnWaa3Uo
sxhvSQy1JDm5MII97o1KQUtJ0wWWi+RMwkIZzC5bwIsDizo5FeJU4lzZkPVBviAaSQNZPYrXEa59
BgZ23QwTfBI7LCvKFwzIUmYBFLS06gcl3/WNBBbq8sGefsoFxhNEgS+XdLxk/WB37TVknz4GQMsF
rRrbJ5nIcNKHAedPj7AqzWYkDlVdRFA2FkZACy9qv8/OcwiIOy1dIF/stwJr3HlTNyyB3HSqqHiS
45v87v10thVBcG6AhKaM0CDZHbahOLIjGfGXOx+1P9GbKZ1oSnqTKvWXosxzSUtwt9YeA63BTruw
U5Vv51VJt0Ht3Zq3BZO4qXxA9wSw5BPR0I9BFgRp/ZpyW/ow6h45W9qF1fPszcTaQO4KAOa5aar4
RiixAYFQEopnK8rnP+jtn8tuTPZQP9WzoF3Py+0Qj/YHdr4isd7RRy6/nEfh0ODS/eqRhEc9Cluw
7faMn01+Pp+Ndjlrp2KU08gcyDmrtll5Je5kgP2EOIVQ7TWLcm9v1Cr0cuiOuZhbDzNUA4cE+X6P
wr4vF3Ca8k5oD4gmZLEPtAGPK2OudmjcmdBLOBFnu6NJrsZ5+YNpNHhvaxe+EDt9lUQK1D2TQYLZ
JpPM9FWK0E/BuxOm6wkI+78q7WIJch2Hrw1b7qBBZu1z1V1I8wpFRN53kfsWswe16v23CZi42SZN
KdjUXd1IXqSi/PNAbKH96E2bwsy4kUfiQubE8iXOu4+12c/qOf40zWM5kkXJKRTyS9/6/t8PQe99
tScC7AS83ByN42Y7yIgHeSsvcHWmhnRedwjhMZg28Gr4CVaytyMaZ2p7b7za/cg60Gno/WUH756B
tl2xs+Ec0GWQ8AZhoNHA8Hu1d26Q1B9ZLHp1prci3hHojuqbU8yPiF/fuqhsYJPQZo2JAGvMRYMj
NYmYDaptshnjQLw9tGQ+9YReKlml1tvQ3EGjGUszoMTbd6vis9LMELbVXY2CXoZ/t8ztF9Jt4vOb
OUAJ4cu0EPFQd3GJre5jPNbwdOOfRKFLTCOCCn6DShRFZP8w2KJPo6s8zzSHTbOxJIbksWQRy//9
NULmQ5w1nZSrMaRZIgHFPw9h2UhkMTF9zT/LNT169z/60K7hNrYItFq7eq8yqnRaAO4SZgwehGgd
TS1gnY92G3XVncWPcDYDO4/gfPZtFXnUdNak1I5TbP50JIYfVgqXfox+90c1HFmac0i5s6NDaJPD
UVuy72HNQKOEJYzF3FiahZFuGkLm4bvslkzkcspbqdWguMpKSp+eCbo0HjuhLbCuZXgyom5/PXBX
7FtRi03YB2soyv/fZ1viNeBAzgmrwPN/QClOhE1ZL4xB189kpuHXHR1VI2knUkJHhtBzSL9XK62J
sn9+WwaHGX92cMoHXMR7Gsmj9JAKckFEHakSGpCScY0Umk2SMb4Fom208+WxSJa518iaFAF0ej+V
EICWexXMaOix1Vp4knEfp+mQwERi9sZR4cJ7bj7/9Rfuq2FrnYTQ/vLsCo/ViuoWIChRShmmTAsu
DGQHKSRuHqjgmOPDj/AZnm1WBN+8E3vYPYCtrrKSEFCnnfUUUFO8zC9n/89c1R8PkFocXKqE+fed
E/Jr2MFWeEcV4DoT1G+JOMihJMrkYXy9f+myZem5fBGecRxGq/M9CDoWjcP4sCANwwVyiw/Ybrm8
NhsWTqFEvUbWHtL23nXphWNQtCPYn4/1cROne6+k2NancvFKnxGsDjQr6xUscs1FlRL54bJ5C3am
89vSfdM23X+dLFTVjDLKZHk9AeW+cZW7ziFnrOEa3Yfhffy8hGXGlVId39BiMA6PeGtYZOCAOnE6
Ch8+xMxzW4Au+ZfjM6yoNMH65nNnHiQB5zP1QJksaZjtPvzCMfMfqmfcLRrVDWlBXTyelP7IY8xv
BTMasjKLlqOggtPIa385yauHu2sM5cK6/GVXlujAknx+4q2QzDiS9wTpPL0/OxIMhGZu3NLtb8yi
OSkCAXJEYgBemDS9DziJNd4HrWE85hWuOlFEe/fgZ1Ci2pVkQm14/DZYP03j3FUEQMdS5Rpp3yYm
Krk+XogAcAeRHMkiOJyllyOvA4FlpL5YB7YqMPWN/Uj2LYniyCAlgmF1kFzVRyOdCr/WMvUCyUN8
uk90X77/9eYFi1BLTkp/3SocEcR90ne/76dJp1DuMRGdlsHHeL1D0ClZAhZr4jlk4CWU9FdhX9S7
tArr8e/HJ3k6h6vv016W4mnWSyo8sagTxw0s6wbmInJyBt6ia3ulFrzNVDrUnZSjGlW9re+NRkP8
AaEEaVY33idZ04dtIMduedygloXp5V0Tt+ayddixoOLiaaS4AJinXpqEsZnK6+d99E3ScFg4X5Tx
Y5ANQCCZAidiJmJ1l/oSmGLMTVqD66B1EsatYXioNqazqW+vJGfchgHntTH5X7n58WvyIXJqj52N
dSeKykYX0rEaf1XlPkLgwHs5rsVbVKK/o+O0G2H3DG+DhP+OBpw2G1L06FxhAl5r1YPGe08HyR5Y
1GdM274gZnQSNsLsHK+vNWgQSi1uIgZ0M5Ey3hpQc8NrDo+pGk06uTPcr7AYuGM0H/RrghPlU97I
nIgR+q6+OFSnCh/PpGTj1Fx86BqgQQJj6ErD89tu+lS767/o8k/9FOGTuMOQrZQCGQrJSd3qkpTV
ZjN8Xfk2Sg9zPVKjnqDY8uwCnBUFY7lpp3E+wnYH/5AMak2iZ6p8o9c9gHOFhKMlrxgBuOpBrolG
aOlLsQXMnbLgHrdfAhTrFfOm0I8fTYTN2zUt0e3YN2G9vBYIdfAKBozOMn5j9SSPIsC0HhLL84Kl
t7wPG08KcOIhECE8zeOz/xv41Cx1wIVchduVii/w3d5G8QdmZiW4Qj2K4XSSuGuXC4ylqKXEpWqf
L7tzfbU4RFMN3cmv2cYhfJy97SXSJcjt6QfO0SD3CM2fVJlReWau7FuJEbXcqgZby5/7mS3hGucq
nA/LEmpQyd8dv0yDLfjlDYQMzqQcg47Gr4aLZZQeKNWUMaE8hmMbgoRUpUGl0zSEA3wQKWybyCI8
CEq18VopqPnxeoIKx2V98hPW2qt3po+XtzTccS+lsM7GuLBQW8smtAktRfuUmsTgkEpAWsmbqQPp
bJkA7Fsic1e3FhEKK1VNLaHxtylhMOu5fqXh0eIFW9eX/cwK6hhKqfXz2Tf0ibu0RW4uTw5SLTaf
NdKJRfaD8pfqTmCqYxd2Mjecsq+XW1RKNubWg1nhobxmWXshHDHmlXKem1ezRRKddJSMk+T9G6G0
Ay+mzlOATEPiGF73Usdc6nKVG/6CzbwrLBQKa6Tm3SIhlKlbpgGWKpb/BGqTGbRrAs+sP3ujYvMV
lHk1IlYmdE/eJLHEmFzViDXGaQU014yKM0ltOSRM1oCvlVKl5uaPjU1EHI45uWKsOXYjDEAoJewC
1thLxiEiOQSnpIIEIwAyFu4wGayq3mdbL4yjBbSQfFWvj5XDgSaIIRN2XajxnAJHlZfxtbhCuAbF
X8oMVbCPICyQupznV1YM0ZyHYeTjdti45FvKIS05u2ARQoZbE2fjFCI4A/hCMJY6milW7vF/ok50
0bA1TSbFICUh79hjGn9IE2Oetps3oEhjDuE3UPUF8BijV1VNcrsGwOxWbcEczmFduawCknJr/EDA
PGDo3Hj41N25Pu2MgDbUpIvGQbhw6NaFV8nzlHvOC9h8g7E0yLRK1Q7Qd7xkgv5UsmhYP1nmLlq+
OhJPtmEhKGfO0kBUgN40KelkyJeLTk2NHHSDmJBMuLlyksnV5LOAM8N5Zi+hok2/j5gq9B7BIRae
Ox0aOpVFmCYw+HqkMAAhYf85cjnTAF0xw+P9t76jOkhTJvxb5s9hn9oXIry0fJTAJXt5L/GtEXTa
ghhB3Y4OvO7O28z4n5pl88dNPcPM//j6hBpo/EE7wVidycqKkr9op23V+zlXscv7gnOJqLfwqURC
p2HiZL148DKgPwXPxJp62pfQriiAoyo/Mmlxsrg59Qv+8vH/S2mTELI+prQBy/EX5wAl6/wfwOF+
l6r6KLP1Eo8gl4W6v380EjsDAfnLbpvI95Z/Pd0eku+Yyh+m8SpKw/DN3Tt0prnpI9po+ZbqR6QO
WV7rE60UcnrVpUQYRrGbtSXXW084yfhQDNZi9bYZpK9Wp7I6WuRUWOpUhspLb3V/INUFmGhwBHp8
DgQcYaSHUD5RT8tMsskpuB3k0H4s/KJVnvQzPAotdFK9kdwzlT1N5GtRWAr9wR0agVxg2NvP5b2c
kJoJPlOLrctGadMF6OZHxL7h0E3FJK9fR4Laoo1ZZHcK61TnP2f3QbCsXqmB8FuPNj6PBTT/9zze
RrDsUhKQw+xO1QqzYUHbkX7lR0fQgSSSyfPCTJmox9Btzc4Cg2176qx5hVIwaLlxDH5sgnsfnGns
M84iARjQekj3hNwdbNuQ2Xz/mdyWeDQ7ad6p0QKRoBICQ4iLAYg0/StJcfWDzec1HW9daKWwyRXk
Cjr+PT88AF0lakhYab1HTXo8j1GAYN25+UfAcXjtCJAcK4gv/DJhLoiXZScP7uPaX8QHqZtwzSbv
/Zr2fDC0xdoXzjXIoCQXPl1hISOe6BIogbd95tXXxuGwgWvcuYj5avaCqpr2sjOV6hqK8X/Z347V
AFgo91mAppgAM1b3NnenKMoqk7F02Av2SyuZ3DvmC7DpJRe2dbAHLHHGfQ6NMXq/Wuc4FL2mlbr+
1PB/L67xF5RHk/VQXWAQ1mZtVb+VkGDZF0biXVaskqttn4mhszEt6RsHcRagS5WxmY576WlKv7A3
PEwpLIASsZ6jdVrK592yf0B1FNFZub2BWWdjH3+1tW7YyzLmxt8JyiYDrBfvLlK7EMCLMKiirZCm
1P0QVzU+WvnADtWGKwOW5xA1jr7/hLYOvHdHobufnYsQ/vTwPFZH85Lm+cm1tnwhZxSGTX18i8wF
zqkmdl8xQjtV0BsAJ3hi4nSREaKnkIUo+vkSpBZjQKEZOg3bIjB0WqRaVuBGiilzQkzvlpegv/tW
nm56hixN1CpKoEex2pGA+6W52bG8eOu6BW3RMBepFpl+FK1IXwIVG1ivAERPVvYd58uANHbSOe7M
oEFRxNXFiINYk2+ESE3qijy4DWThiWAD2aIZ2Km2NSWreacxPHSCbNu1zb3jevXWuJIPEax0bkRs
RH58cVAYJ0ZKVWqQD4UoU7wmryd6HtnNHmj+nbrGkhQhB1utf/ZpoAFzwQf2Ene2/yKarCtybDBb
ASckuJOC6PlNEhe/Mye5CRVCMMpg5orTl+OL8T0c9TlBJNjb1vlRva2Rdrfi2JVwOOjmpVJEdkda
VjzXcuXbo3skSH53XvERRhlzKFJlwsfGBqXhVNO+WN/xb2ifmvM8mrS+MbduXaipCDFcTLXEbw0v
O9tjHLn0pnys6E91OMyXjV0BczBjc4Kq9/H/XWsznj5JJsTv7qBDG/8j3T5cuyCeCruCTrowA5Rw
osKn/szu3KHDvXBvJDMvjsX3lx9ve5IarvJlqHjCZi+VFQS4w27eG5zX+qCA+LdZjIthQI7QVqG/
bRIFRvCG7k/XCLy68nZTBr4p+V876tK1c7Rke9iAYbC2BILGLyAQoUeWuzt2QS7D9oZ58o4J7h5q
+VlZ8tPkpgpc0piFIiI/i7fmeRRg7ScK2DwXKaJjK/yGnuRQtf4moJVWFl1jdrbq2aO+Beaxw0s/
X88zItwR8l4fUT376ZzQTczsASaKi6SFPVapy3dz5Xy02RuGNrrE6440bCmdXz6vuXzza9VoK10Z
U4E08AS45WdKFcVUPA1Oj1elfrtuKY71EDSnX0qbuM7JpI8pqbxVZqLlycx7EoBDk4YuLb6JVXER
VBsNDpRqLdACB4yDck3Sl58tQdf8ak4CyyjEzOMmQsav8elCIXXFS5a9AJz7eLLu3p84a6uHP4ip
+AjEUoEZxpQ2kFyLv/BHMM+7SjjhBG0kKEwyAfdvbaZ9oJX0QgaF6e5zVKpBT8hhCS7UA7vd+l1z
LPosBJKgebyLxiyaOVXWcYtjOsVs9847H/gAxTDmXvjnoeXX/+xYsPSjj0bJI5Ip2jQyAcFX/q0A
WwudyXjaxSqPtgaDKACSFKVIhh5X7q9Ier0jG6A0Me0S2vubQkAqryd0+mE3qQ1yBoYAh05ZKh1B
qGWHLPOMV18VS3tDjkPHGExfvmqWBwn3dS3x6YWVeyvdHLUyrUXGGgd9+5gbnLZUA99xjby+LKhF
usIuFk/L73TIvKjCtiDAUApyeJODZhXssaHZpgSVwhXPZtsKdpfhfGaFfRyy1Ok5owwT0wN4c32K
AI2reSUOhxWge12tUQMF8rm7MJfFjZ9/RJuQX8ojs2zmK9MNVbNDsKrGMviGkU+F/PWL06ucQvZp
b5KeciaN0ZQt3HrN5Ko5+6JQArzy6PSHNUSx1vdqY+tDaXSyMvEhmAisI+9UHJZ9kYNdwvfGpzmj
NfDOHLy7zCxxIaMPi9Bf7ysy5dPOkSsVgCGIBXLUhiI+XsDYbnubpygvLFAgBJW9QEoit4MniHP0
8hJb3OH5w+xe0cdcVCqubC+xmlFOQpaQbbsUEzZR5Zi5DiznhEj6sujyoFfr9MO0aShFEN/ysZbh
L5vh5bOpt9IW9a85dD+u/boSDkNqPwUSZjHDUjP5lwDVr/s3PHoa4fSWveUL3dQyd0X1hZr41z0I
nO/gdd/Wz2TxqcIMu8bMf9n1d8wABsKaBwUppJUkhDSHmIUd294d67U/oyQri1HScCBCPa1umG/0
mmGucuo4z56QFPDQ8QB+jUiPYXVKNh4oHO0bma56vqfSh0taLItZihfvFucx0rNdS871ednTnUOd
qrVWr+r8LjHkIkYLgoRvim2npGek9f3vgwvIS0u+gFLKCnSGd4HnJ0shHZg3U0kLBIm1avJkpDJr
sgglj0uxTx5Ovk90yJK/Trgr/8sqvCYyVqUH3sxTwyRsaHstCPIdqs5/ORh9uQBj7U5Q1DM23fCj
idySoC9LxWdMPrts/a4WYLxmkZ27jPjG2mYpt9/vzlXS4/S0DoE4Qm6kLxPNTt2aFpY/ifP4Mak0
xqrnHmmXwvEqNd2E+511Cs6YlCEF766n9QbK8EXhNHAM4ET+iFxkThStR/IlwIeR6ZdwEtI+KcMx
X5M0wPWXkUd7hO09ZHp10RayWE9OEXP2WAAH/Tg6R6wlaPAX0xP0NjP6o4t8SaZ9WHmpZz5ONljd
TSN+fnj9+cq+YEkjdqdhrErkzvv9QO8HqcY0do5AuzhXL12n1dn4Xl41pn/rdOHrtpAUwQYt3Mqs
204jsX8GXd7fdRJOKN9nsvqrEtKyebh7xE2QY807W6s3po3N8jKMJjZmjLPTFHFoSYUBz4n3JhVr
lmLOJoGlyA+c8D0z2vAtrOCeirZovllu+rBg9rkfkjJ0RgwTN9UJ3n2yU+nANHSjHrgiFSw7+YmW
Z8bCCzll9izeEyljJ/hB1l9kA4i5EQoJHO3Q3RwvZL+XNqLP2+Mxk49j6APm1TYiwz+HzenJQTGQ
iMnxmWYrHXNA0he8R3l9SuBQGOgm6j7OLQM4/2ob9wlPgGQZdrf6X9DgGAN8n90a7lvNcEoViKxM
PUx4onl6flaYwl5zN1OjI+d9hry22szikYYZX3Fm6eBPhAQyWx5G/u1ii9cBIOOE/Q7tKNjtgN8d
TAjKifUzZDh7MgkVxEamHORTb+W9YsGtqHsRjWPPOh4HTk6dGWPDISXOdkQcyLLkaGlYziC4WZ4u
B9DHM7eWwv6i6tM8LUkVwwgJ+czMzZyvoqfwlDa27oIGFpXGV6yBKng99d9LO9NKZTlx8R4mr2Kd
EnXVNuyk26zcaRTY5dkyPyYy4eaNWhKcMJq3FdN6f0017SotyKhPG1q/ZLvtigPQuWsghSpdYkIJ
gRZaLiKkEIV8YMcxlmjk0d9T/wYmtVcpHl/MDrXNL4w8RRIw+OjHIYTIPcUBs212hzevzzHtv0xT
nMuHlCYAH1Y2xVlEM1IXCGy1HrdJlhmoG7c4vO113L3bhWc8CLxfutXa6kBBVSONkJmisF++qgUl
HqVGmYRMrCEwR3ndHSlEdBRWiI2vaK2wtwARco+HiH9jtUyFb4F62CXS+3siN+cOR48gk7qBrV9n
J9PJGFL9RSD4+N6+wD++BT4nVUFEba/68QjXHF7rU170SIdUITSTc/YPG29IMR2jEN9fmW3O4kKY
DEkAh064iYN4H/jiZbHJT44ZiPX9wU6kuCzhPVhE8BdWYOU+86M2/jfigT+0vLJabv6xpeUZ05Eb
BIdh/8uXZvhq8+wIU3LnxlRgz1bBATMsJQAPjfhWGec/iWb+Xl1G/RUbbscX056heNumc+QmbTCC
RY3Mv7eRmCp2eL6IdzJIDovSuOonY2stJQ7u8GvuqtBP8YQNXAySVv74muKmTeFB2O62X8JLdjOs
wioegmUqTE77xiueyimFFGWP4Xt9fL7/SNX6m7WrPrc8T9z+xp8RT03Ei7wKZd/NuUJWx5R02rwB
032Ey4TMhfMSHNiWJ9uVE/xUVyUn4ve8O16JOnA5L38I0jyVMLH6dEbfN4N2z6P9hwHBQXee6g+s
Gzn1o0N1femRazyN5PeZICHJPIvsNpmxwkbGPmWAETErYNq0nXmviwAwqEYToO3lj8CdlxfIkh25
RpcWjLJpGzSXrNxkG4vTutBiSLlXnQ5+4XjiohTgRUAPP9f/pgLSJnENQsn9zQ5/Ajb0K8Xl9ldi
Wun3vH13JkR+lxUYOBIjzUMacTuEoAShiShCcUNsWdeRXIBzvM2pGNyNpMQFoi8KoX0OBRPfchjj
72zeoWL9DRqHu10vx7HjNXBNp/nmRTQ5YUT8uSNnZjEqHmiYoJbVWD5nZLMBhyziynt+usq0KlXs
zuXSuow7820RxRl0xKqOW8eInt4b+hiWjYnWbjQ7jCh4qJ9w2AYn3hVwG7EEpn6EkfsVo8CmQZdz
pC2Ksne4YJ2VXFxBWb21dzBYDIPnMlyk72BPGkvYaHGMM+tBULF3brtz0C4owwDvE9MpvwJtxDcB
F7Cv6L5bYGO9nXYavocjvl4OXI4Hsh+qPysFhVn++JiQWk7ONiwltouB5wTpz5lgmGjIZFi1JU/h
n7Dfanqt0wxDWZpTVip3L8Hxj90FgOlF6ZVZ1SxZHAdI/6CsHp2+zgSPZskm2Nu7BmX3fI8WKpQY
iO7YTqk8ou6P8sDwL/USUBxx0oRfuGZs0SotPTXUlFKluqNaUz1klpZlsQ+6RFy8KaSYvdH06sQz
eCwzaa1kCAdc4vjJrb8+Zp2Z4ILSggpe/TobPV53F8O7ObEZKFHvLCGSoWqtz0sXCnxai0H3dUmK
mqHeUivDBREvT9teGsp40CnwuqC2vRNhS5gVNWm2Dncf3PfI6DKk9T3dUq8WWcVqkQu3VLlBTEEE
sy2Dr46DVnmMiJkINxWWanvhyKeoCOPXo2V3wnxPmC6b1Ipvd+frbLMBqcD8u1isu5EuFc2jk4E1
GFu8iVPGjVVfqWwCgC5eKPNMmNL/Xt/1NO5HVR2ZIVEeaJtOKfvS3l5EGECz0suHzXOec6HhfDwo
RliQ1gB8P+j5A4VH2BiENtYEUzcPZiy947OihcQTGy6MEpackrePWtK2J4NB4jF9PTsUgLez/GEq
1VplQzz8aykE8C9cs8U6eqWEUYycEzXpl3YHD1pB9SKXdNFoyUGRUX8q29gLBnRo9W4jSasy1NSq
rbI8G+uX0ZRk37SRpyylmjQW1on25Fv0HqwrHTe8M3ZSgcBAGAiCUrE99S+pdcHYdGSeUWz+3Xk7
2H/sv9MB9pNYOLrN3ElWbuzfZ8WifTFy2qmpsaOyisgnJGw6Q405VLKari3gQZ+XglKTrqGInbz8
9Bz+ap+l4XpKttMLvPNC/uEzbpLgKYYGSe4zlrzU51ykaYT/NS3hmrQZB6wv0ORpsLeXeq501mU3
D9pfo2us/C9aoncmSEz1EsHsoBgwRtTUi2pd+Zk3ABusN3j3QthCVYpC88qobFWAp0wxoaTpKWYp
oJ6Bcr5Bscj3DjGG+gR58lwCAqpcnuz+5uGn665otUlx6kxaTsasRFkO+mRyGmsPH1yxl44d/14D
Pn468n3VY5Ax4YhSCVDa9G273rrBdGyRg9rxqsmPUD7l4LXE8gw/qB9zZJu4n18RcTleNywqrtwd
iM1RJ44rESUGnCE5u0lbOIM+jgoM50jbNc+xkj3qc0cTx6+nZqOS/9B8RjsNCgvzleYrZEslbGNI
Cbb/GY9zhUWXrIvAGCTmcZCiuowPYM7ocP0ZQXPIL/78ntzmepcfJIomQ4gxT0FLnyaKfK4aaEPT
zrVpQ4axXMJ8ACtrSHfhpNfyGdkV0TIVD9iwcd/MysO+QdUK/FthfC2zwNrB8BIob5sBPs5YJG67
GQLZMbE1t5akgI3Uyx2ur1d1QMdvhOz8KCr0KbY//MR88B+REm/Q7EEdVXvfzb+AqyoqjtD1T1t0
aUEu8xEncbeff6kJnPzq7JfRRNkQYF7/6SdUQdpeR1S8ddF50SO9WKXLfGx91PXitCc9kRH1skKq
5zs0o999p/bSzgWgsUQLyAnH0aTlTUSzsNxdypfC57axJd2Nm08niktmfSLn6AYSH5p4jSy2KhRy
z4MXWh12LkHNlp/VWDrHXx3yzTnJrpfpKiu6MMWcDWgeVrkCq07WL1XnaseLoGddKeFrdZyW/woo
BChHlYPOdQ7FJ9Y2F/HFTh5UFx3JXfMOplGJKpTI8dcyrATtE4pWYD0MG3rDPCpvm99QXgE3iocP
jVtkDiDH+Gm91cNeT9bF5sTjfhFGGd+Ed4tooJCEWrcF7nmsRu+dB6z1cfqjbE1XWr5Epc7pDE7F
yDzuu4kMmDyqNYmqnPdwUaA2B+3Iqqqve60jLo9KXfiSQsnYDsmbc4TpVibYmilnAr8+pDsoBPgU
AcaRgZW/2ALOf2A4zuZZzMZ54040mDcYD3RMdZgsDPBWRFE+Adj/lC/xi+NfofrxgSSbFjUNEokJ
QhaarS0QhXrlXr0Uw2yXeaPI9EhMl/ExfrVK5xLiWnIwvm17TauIt+SsF7p8uHQQYEap+nbnk0B6
8HdJhXRi0gieAAB4ccOH8wA4czBPM8fT6nMuTmHvs++tJlE87uVwUsMMXDYFGB8VCM5bdLXI+a9f
i8OMLypMFoPEutQZ/afsVRnPRMiw37DHKfZwojLmA63q+zncv1KOjZi3Z6tZ3fAxcRUcToK4gc/X
DpONTLGDAaAGbDWwyKoSu1cuoh/I2UMg4gBXHyLnsKuJuiyIlhG5bySTJhgNu2k5bx6KCh00/SqL
UruMWb7apS4+s1GkKjCMgC1buZJ3rF8OToG7Aj8kkio0kSGmrXVLvJQ52iJKidFFXhROBR9Txxhg
iuXPBdhlR0M0QKjMlDNxatZclLExRg9HGA9A53wI3DzLYLpeP8tXt0tUf6W6acUCAwGjYuB6dh+V
iVspoD+too0jFeGI5mbdxky7dTCCOf4JodNAlgNAZBKPrbEN/+LXbCrIB1WkToNtz4yeA2j6f/r2
a9peO9DiwGyPQC8/LJMc2RnOczMuJxFmDX1yOmQxCqIOfA5TDBXYb2cGlZSfj0wgBCXjMNDPwTHf
VTDWKcrIGPgisUL+/7L0SE/vOvS9GiAft84QDnYKykbsNOmvf1SzwnVEbaLiHxlWiDjYbi5dGk3f
tvBQFThsWVURAT5TUh4a0zkpFsiS3LTB+pyv1TnUGvA17yfIGE8o8wubjN+Biuvbtj768wH8+Jxy
vFDoaD9BcAlrr2Ki9nlKUjsFZCfgmBY1sluXk+1EX8QOFJqcvgiaRRW4btMECaZmeC7YpxJ2p8Q4
wDC52j9FAh9nTMIHVpt2vnhPqVQWaMOOTJ3ddbCuEyrm3eouMq+xUwr7IhDKLnJ+GWrp1mlzp4cZ
YY/eHrOyBX4JUJrw8nfscAQ22ZPjsTo6RNKiE5T6HtyWYU2etB7/gdiPMVlHtkUkVTB8tl1d03oJ
Z7JL48my3SIeggDMDHyhqNU2XmjAAsKaI/YXUj1NsZoXqeJOKJfKUd682Ju9V9Q2Hxm/N3r+mxc5
jsCuU/bKzFFobqWznTnixsXU/kXE2XevyezPHwcTGbR4R9QmgYwiEodNZTUpMOO4ENau7G48dFqc
al243wUAyaerDUSOFUHnq8wYzLkOHAi1HHL7HRFiDrnp0O7awdCsRKr9rOnitb18+MkSSXaaj7gT
S/eV50oBul8jvQXdn30Rgm7vyExKCoS5NPEupIgu7AErisO6eOf2F97JTEy0WHVqSzrujoMqxn6s
Kw5jn6aCZSxQaUmyBb7SYM9Le6bogiMgLKKAXUhHfLyPIAhsjtgZ3dEwGcrlRKE1CJarWud+sEMP
UdfWMFWmWOfFoH5kYrnohuCQtkzztR7QGYsuBbIKzpRRWgfWMVNFCUvi2PZuIRxPqccJTu4wsB8R
ZEtU9H+48FrzXRt/C0Ig3vo23vKQ9oFPnR1pOlcjBmyjxlovMy6WmRILxBZjgGS32wIv7Y4tBhgs
NubwZf8d8nPlGPOFnO76W0Jl2JJuuMeZIQZdrtU7L23NPAsgmAYOyxpRELIP2okcs5N/tt5TujfQ
sZHlRcQhHnLXrRfe+auk542l7qCi7IZc6lBnAUxfVh9HyIko1VUrQzi7l4y/8Dc9knYNjqVm0jhK
5rebY+jLb+Q4ITHIY2MbNHlIyWVoqder5RCboGSg5auM5Pn8FyOLTEVTwtdQ346qWppcdiXMnbl/
XGTs9je1pjetXhOJ2qJkQ2alFtnkI8w4NiSKmP9jIg/jQaXIFWGMfdFrF7Hs68YQN5CBy6iacg9Y
D8fk8ycAVzC6XljQqNch8tkXOcwYwIu9jZZospQdq8vj6KnJVz6M3IYCChm/jF2Uzw53hCV1IiCd
cse1kwp/QNGH5vLVa1EwxfOleKxXLryyhwruoFAf4kEVhfQ8t9pjvZWZbnsJXyV+nmnP8LSlmhey
B33DrE5NOf3ufsF3xv508ArU//LR3p4nLMVLhLIFOZKgqNg9MBb3FFzpX/p4kTEBBwC+j34GzdzH
ID7fvEBCJdPaMJDb3WzF5wYNia57NF7pcLzkoSIZ2KcP7orf7MvGbdvAeV8VcvATZOyFhp+kcNYK
1gM7BUa/GVbJin1R+zq18ocf9V5zzGTFywx1HeH35SYuNdEz6dM39exAvfgrKte6ssjukNkvKqHX
zUMpBoWqdmv5qKrq9A+mu1r5n2rYWnWKihLXeEncufw1xskpJNI47nlJonc9qNQzyXX4K1tp7TCW
5Vk3CJZHvrcrd8/ZsH4ZZkDOyoZxhIzLFBWblnRRh+t4fFJvez/yp5bdh2OmFZMeIeEsfq7Jl5Zw
EStXUgLs9r1NJf3Ne9aZRsvN4RvN8b1aLVJBhUvsRbhvpCF54F90WUFWC5whLldOMq2OVOZR9s0p
/wHlavoW3yGiHeNhMo8v0DBPwTbjr2xCbc4c6Ka/DKP6Gh/2Z4iOK17tGXCS3zninbxe2vXOfaCs
iDRYg5bmuX81oJESSqnnv9pRbHa+vsHXKEuDgKELbrYRacYzYaUAUygHWMhz3Xa6pQBsztvzrGH8
CDQ07/FIbwTB3iRnMRUkm4v/8mubRz4eMWDlnHlVgnJO1nA6EoJfL6tElZbTaaSpA5j6Vstlmwu1
DE33G/FoUPXTc0KGEONRZrh4UrrkX6KhYinBUFEJcPQB9k12SxbZZxMXLS0CS1nP3OWEkofa62A/
yUP27Yfid54LL2hyVipardSeUAurJdEoSp3jBTabrq2PruMbD1ztFTZxS6Ob/srmFveOv2DRnh5h
JPT0eZT9CwPe6UQquGfaTeGr1X0iYpbgsDJUKrw0I1mJWrpLigGtgBns41tYVAkpv9uiUvQLAlhh
dLy+q33Ltuj/ciPWHmy+CoPmNTJJNhxdhtG63YuO39enmi9RUGWTUdBkz+YwImxg82MwJPTC0rAT
ZYNsAdBfLGykzxCW0irHMs8YKeYxDUU/5x3+E9lnLZu4RP+4nlxVIghRBh/ydRTUrekWwefHi2Kl
FmsvRcDfnmEShWyJFo5l4NYO3gsKIr+9djFE8gNq8Sa0+vly5wn6PXnfXpTKzn7B9FVIZgUWJ05U
+GZiSfUiFUFn+T8hSLAffmMphQOMD97glKgaWXKZoSna8BhiOzrheN4nz6Cty/7SNpUtQdD9PYAc
umoT2ZCDGDCBs24cRWkE6q9RzuONGPZwhBT1oRNn7ssL7WwObcFQkPfwkCeyr0cdJVJE9MRqaeJr
YgmmlIdF6JhL8MYyTeTKX+i05ktqku/FEIf6gXUjPeZispZg851YEKzyB3WgekE9o7DQqatmHC3t
+oW/dyZRkGtF8lRkNt/Huw4TB72Jfc9gKjen1KXSqgrMCRlZp95OTdOU2cQcvyWhOCV0FLHIymj8
7+2Pcb/tT9By3rCbtmI+9s1/ze9eulVVH+r+/bIysz7UJNEnzeAd1zkLuV5mMAR29Y8qoVfSWid0
iKrDAxLaI/8mbjKbAkEmSIl2+ouo6sx8y8QgI3RKnOwM3hx3P7JyLulbuCFGEhMXkZMzlWsbKGAN
7hdd1/Bd5W4JrGXdwaUR9DpHCq1i60CE/yIuh5QWA4OuP2A7PgmZV7O+vo4LoL2jU+K58/o5A+t4
mUWytOswAUcMhhxWjVLB1l2wl9kxZlB6zokccwQ0ZVj2PFDofVgOX5NJxGuO1SYRmvbsoWxe1cOh
cSgdntMs+Xp2Uo//yQY+Zl3jK0DHiz3+VNeLnWBxY5Ytjdbtcgzg3MPVANb49q8rX+zryQsLStDv
Y3qkfkeCeB95U5NwNPGBZzuwEBjSPQYBOa0q9xATqqpvW1XvHpO+wkpjuBSzMcXU8S5QvZsvD1cE
ioT10+RhvAs7L4vXxJpSUl0xaRhLFbVI6b6wavxE28QQ+UItD4MtSo/06daYa7B9hV/fgeoFIFO7
cLBD2y+DqvbgjZIVsVvo9wPa3G+6usSjEmx1cKhQq31SwX5fEwNbqLgkAYeKrtFfjmHeBf6cfN7s
ADxAYlSPTDkvAj/HR+Egh25rNu/j0E62gnc7kgJiWqzbifp46m6frzqB5skF5EuCgh+FqusDloJY
K39X7S1zurh2SCrT73Jyn9j9xSQ/3lXIr9NukxICNMK+/brTAdeTR930oIJtDG5BaZAASoQ09e2I
3ymqrUhpePyOpHC8+hTHIWpQoUQmeX6opfuAwlDXtlhJPhAWSJJu0cKIHl0oaMqJ3yxEIg3at29m
gatX0/jGC7uFviiu4qQ9wzMHGwULWuLq8QxWRHNGQkChMzfJ1Jk66QTVkHBztFGaa28cbrUMUXpT
P3iGtPhCuvKfsj1S84sP+nWGe4nqtIpx6AqWhz7+MJs3KthHhyj9F3TGi4pY/MJ+6og16fvx57ly
Kz7KB0OmkCZ9UAJnyECJ3n6dpJ/P81aJiHuSFNnK1EpFrqr4nCUEJAFo8ZG/6ufRwzrlRmHZBOiL
2E2xlMolbz8/nqG7+ThxdqRXNlt4Aqu0T3kU8PXrm54JonV3JvLWrxB+jtQC3MTyR/IZqMCxGO7c
+nWQd+wZvLgpHwBVNFZmeJXZUeDbQlY8WXSMhcl6tGchfZEsCurykZX++nV1rISYV+I18+tYmxeX
7cP/Plsrm/iDowqgukna05X3EjB1aCgbs3upAehdBIvO1sE7kSB4W7PT314LNyV0DoJmyw9La6qJ
WQ9rZoTs3QXR9AFK/WFwhQ0Ggs5syHDADpgZH6cNtzMYHimnSxuTtmaaJGL+gnxEkiT0k/6m7iYN
Bpqdc9ZJme5BCSN6oypHPPQoPz//HQdNwUbjAUqZ5+h/1QcNhc/eKSr7HTYIeFHsWUU1wEZrO2qt
WcogpaGnxz2n5GrBXOCH0q7hm9AGwBQMNxPdITYjeEc0dm9JqRy9IKKt0zX3RDH4Gz1BEhl3xR4P
LrGhn4NsCEwRoO+cSHL22rNM4SfKv8NrCuun7xDZ1aJdUZCaGg6l+5452Il57XyxnhWfJnYX148k
w9kTs6FbIN0YCyFevfXTlXx8cKfxtSQnUL0Kk/hK/7iO3kYIyWaxNbk1/jsCDxDOuqvQg7bznMrM
MfBOIYycOoObaki6oyLteC/RS8JRwyxv+za47I+wPx2ha8INX8HEp909i3lkY7cQ3eW8tgClqTMO
6DNTrnHfXfZ5odarMIZCMNdjxMGhteJcQtRb1/yMIdGaQbkrlvrijleNIe/Cs45yMwCGD+X7m9GZ
kEjqD6hdCyV23oPQ7Kl4hDhWTzBFT068YaSoG7RR+vQ1o2iNOSLgrL05k3q1a1MReaUpgzt7+Mve
8dCqSnhdzyB27aHTmaRXsKWLKxyJVG+Xdd3DEEy3co0v0QtV0LJqdO+0Kg4w7eHDQJXk2tuald6n
vM42B81C44pU8xCxDoESgqLLUE+IKpqa48tQbDDbnqs0ATsdO+fspoOa0kIefo0JEO5DaKYGs3rv
iPxNozuiIqk2k5/vYFaTv9nJCjSOfCzm2W+72gFa+MvLpmXCCTkVN7EsyjZV6e1DsIHyvt4F42bP
ytxbLTDyF/5p0KAapWtTM/TYfWbFmSZmBEltXRBHGpt5zZku0PfqZTa8nn8/QKSm7R4aHSIZjrU9
0XrxHf6ryl6RdHKi7SVhhOOxpePGeMtazkk/GwIo6Qsb3Swxhz1MES3/3fLPkRKTtnFgx5ixK6Ej
OMmQX76hHsj0MCbdhcLaXIcXCs1MG/j4v+MOhapCuNU5xFvCvIqp8ib8bl6JCCuFJU7iFMNv5gsx
Ui4Pa60SjjUSshZ0UjUyPXRM3Sn79M9QjlVP37xJ80IAwdBR3tdo497mNTFzfydJW7aZzN+JYJXI
KdQTai3+j1TBD1/jn8yhJIcx1oevakvbFGOnI5hCCARBAWp5SnR+TdLKcdW1/Se0Op8AYMb4SMl+
vaU+bXmMrrEgcT5e59+JSumrLQZAPo69/kfQNeu4OZdIIsh706IPhv7+YS7I0AkaShiC9S9jbIWc
ZxYVywZGuYX65dy2SDMssfKs5ioGZgQbjn/+i+fBJc43OEbGYWSgpvNrii9+oxRCaHR+gm0DnPr3
ZrSpCWjipydkuMv5sRpqHCt4tT+6TtZJ8pIFOpp5d7GpTUU3jZBKaqG5OOglLGVrUksJXdsLlKmC
j0kd/2YD4KXyFsJWelmxzYYqYXtkvEVF91Z7L8x2wBZomRjxlzqZXTIk/Cp1UTBYWVMbmwIUdO9P
O2ocvAhfN12SqiszTeN2bedFPc9qjtJMNWFYWtGJdQ2MNg3QXabHoNZiLbhNHKZD6cRTrUAjd+re
3kT+2mvimWw8njZKfQVDV595LhW8usI3la87HFHJYZDJNL8aDIVG2LNtHOCfMurBZKTH4kAp8G5u
m+BQ9FQKEnCxtsInXibagU4F27VV88Pkr6cloDjvDOqtsnAUlsYOG2OCI12u+iV4NCxZMFDerwMc
+gBwEJJLjBq9nhj3JcorouvzAsy/DmjKEI/ofEk0WpqxervKBp6En7Wwwc6fGoq9ml7KI58no8bE
ILjTYINE4F5k/PdnHjDvI+1+m8yKXbZL5DJZ4Enoo7/5iv/r1wbs09d18z+O5bI8Tly3VrA4Zz8+
5IrhM9088Yvo5C74rkV4/Jq2bHC4k35uT5f1B3Ju/1mHB3ch1q0cnnh0IkzGgmydb9FZbsSmYkGS
jiYYPnNgyGDykBUQZMQpu6MCoout6anQZV47YWJuK126sWrYQFI7NMjv5IkKm5+FpAhAh7zjy5gU
xS0/ueF9FGYkGo5HfSEF69QIP6PIJLQv5dYdC3rCDb7o6T6Iafh7SpyRdAHNeeWZ3NuWzgG8yASE
COPOx/56AlW+qAyD7zxrM8TmhpMebos08gbEgqjj8NzMH/t8zzKz3Z2R2NUlZodEKnqRlvgtxAQk
kW0SBYKFFVk3D7g30aSL/DZuMUZ+gK1ZLl/0LIJ/5KaBIa1NnYTv7Is5cGOvcrlFlAXIlpGR1VCj
o6463EN95PdSX7z1vQuQJvqp4w+8EWslETL2R+RtR7y0WkSlv2i0ncXvW0aHIuDx7UYahkX9S0rr
URENpz0/KH5U4L7w7iljh9osdZXwD4nNGdy6dLGDW74dHljhD4nNejKgcvC1OCS7Pl6DtocYeTs8
SaU+4HFYHT9wXR8v/9acpQruEmF9PqKC7SMdzWnDSXjMgVoqlPHk75HxZSgHSWyZbEJaeTIOLscs
s/VbQoC9TpoABXr4jiHp1NwY3PRSVmT/k9L/2FOYp9/PSKzCr8QWDlHFu9odI7sh5vE/dp4xcJnl
m8IWwymjKBAQ+OddeY4W1pNJK0dfT4rGo7scw8VFHH/85I4k7FluT3gRPCOLkfkW5Ct96gvQvWT7
0hLRwDirtVWICxZ+JRZK2W4YPyrP2K5z/i8XEaiVg60bX8LYFwCzc7mjKDi9J5BbTVpAs2p3AI48
GnWglzP9GxOCj5PlLX+Pkg9wZjfRXhXqHnQ+Hzcn2Rp8qjRN5G5jg2BmA/qE33fWpeg+3+slooj5
ZKjtS7OehW4YpKqQN7L5elRTh0EtaSnJAX0DcFYgKyeB5JFDkN2EwvygF84wp1fErhYzSzV2YnrA
QxCYr7YJBKhd4QKdGCWesoqMCkbfNIRWHc7Xx9tJee0NR4k0y+XtTQmxHLG2TvNtqgzfMiOYx6vu
c35Ob19o3wV/4z1mvTtWZ438/SrtIPGgpeuDKyMa/V4IaMPujDjZk76Gze/QQeQLa4qrl7wmPKYh
+HW19DQr1N+RuJP530e01E18aFVpNx0Ns3IU+vy0nS4QC4WDlSYgCIePjGTBpBM0MxetpZ8cTzlL
Hy/LEdP/nft3AF5E3sWbTE2uPHgAZwll2kVjUQcrXxDWX9z4DDCc3MXvbMWOUBk5/WotPG1DtOWh
GHG3fPb992R3bAwO4wHYwcEgWMvfXm9D6iPYMhOBJOl8pPZmQoTm23w2b0Oqj2endXXutuhUTq6o
A6Yl4g5IQLgooJHkOABT0qZmIN2Px6ZcqU+lYmn0z9agTdlV/eG8il2ltq4R1OhrqtCMwoetsp0n
gM5VZ7mTHW7UdU9NLsCYDEXan/+of0uTLpyJhEhuloRpXc5CrTLGEdh6jxN6X4GWPr4HLUhTpHic
aBKmoBGeokQW/RyEv7Nfz1CeA+73grr/rbcxoUl+E9xN6Vpp+OF1uNgs9dQDHnBBfR5qskCwrdbF
+PitXwG5VVd6pt+qs/ffylJssilN8RkUN9Y7kAVjq5BsgwD/8s3SwfXbp0qOZUm/F3GpaRnO231I
er81XUQN63lFDWmCT0vWZq0dSYfe7GR7sM+nRMM3Nbf+820P7j+K+Fy+/Dc1Y7/3zJn45fsOUZD9
Xu96uFG5B2TGRVdztefOd0YHO91m79AA19EZdBLawgCo7kK7eldPEl+gIoQuYYQ4XTuZ50eTl45d
fijzd03jGDMrfeIR00N+ckHWK4h+hyhoquqN2bCEkqd1xJwc4CAYFC571XPjddn77FRnMYfnO/gf
0kPCzCTvpMbuqM5Kpq9QndJc8w79xNra6KHhH6DXd2gROmHRBp9zsLYlccUXkhdaWdWODASy9hmP
qmU7vAkhQSmftzcA+y/DCCV3xIDTtBXvHtXbFz0qDmzDdTmOXfK4AI9f9FWCJHE/RpW86e092MJW
AZSRukdzDV/8otiXO4EoPPeA5ZH69TqfkD55ak748aDRSu+53oPaM0AT6b5H3N3ir5Wo9+JpdLBC
lP22emjNIQyEGZMBJQtlIngoWoQFV/FUQPM/IPqjZHfwF02EGqZK9yXVnqkVTuGN4PgMJxCp7Npq
J3FgQC8Hb+HRlhM4XJ4yORgHKxOyhcXB7DmfoMGBkbr2OOfICMEJuf4sXse9+yIWVzdWlBC5HUaK
QroIUDbYgtKpXqf3hb5xDS+2xTQSpbnz8/clxVpH69+ZSoa6UXurHHBs/V8yrdTrxLezAbb0FYo5
4tkYj5nY5JQV40EoJy3MnaPszihtwzsgc/WYJXDsPyQ/I1dgzqd79/baV2m5Hedf6Dc2x18XVFSN
COXU/JFQfd4wfFoPALpTf4QFwmj2AbPPpe7dK+ztmBYa9ev8GV4tRxoIBD2avhPvQY9w9CyX850L
5nwBcZJ3mI+doazAC85E4QbT1YLXm7GNkGXhgNcN44hddT8PL66o+gTXlMvUy8VJzMkIJyihD0K3
J/0eMo0KJGz8rPVAhVmu1HQw/LqEcSjWyxnnYiOdrC+hEQgXwvY+aSDA4rfZifCTvUkHJhzlCBN+
T4Ol4WOSUMigoN4jAaAvFwHDH7ZREUCPcXHmjzYwNBARomiXVYtL5Xwi1+h3PXm2h/Z0DvrAvhsO
MbkRS/NKLNaSTIPApG5MUrBVT39RHrJxdBtlVeRnk6NLVYsixnKSGrPU0kylu0kpOkWnO4lu4ozV
1v0RavIMGHoEkqtJu/5Bmluejm9niwa+Pg+cRTIIsLf5LpdQUhnOrnHJ9mZc6aACy455h1TE+wNY
Pwkdg+l+PzG1aQTM3vxBQpgLe7eovuhloANUY05AnRqubJZANJEMbhDqzc21R4rDLfyIJ/jrOHhY
0zAD8BJJGIgvneWFZVoX2W18ML+D3g5eZhP7Cf6alEnlGJ1RXWZswnHMYRaYTC5okLEyxr7O0KSo
XpkRJoXuUfHwADKdZFIBqzjfaYsEJrIaG0s05lvMIwfBBlL7DS51C0My+oL+DeJ4oyk8n7jH1uN/
2HxftWhrgQouPL6j40hVtV60WSQGMyYKb07Y9zDYVVodHC0pkHpCBmPYaKLZtgflcu04SXt0Wo6K
eFFAciepOMhAgEs6MOfDtIbSvMqRsRgleoC2kuFW45ppiQJ3QgZ/WyRA3uGSz4djbETPJ1lo3B9s
BKapZJKGnVqW4mDwnSvpPKeJ1Jr91JR808u4KNYXT9PjNdPQeFNceKoS1woCFy2Nn0LQpDOU805C
LWYvzoQqPFxTzkw6EnIbF6dhrmBAREUNCx+PBLieGgNM4kLkSc8EsN5Nc3V/1IaTCuE4hzzQjBBo
aE59Q6AuOFjQxzvcyICg1Lb/LsS9HwN9wDkcfhOHxgp89E8W4GSJ/IRz1Kf8eKf3j7jocwkImyLB
3T8cipEs9KDyUWPJF3aBY6zw5yWhP2qCxD3dhPIGH5cxzEV9srhpJCpxfgBQ1nQJPNUhQPmFz+lY
392WfXD23a7WwLW+Jo/jtU5m8DNETFzoGmniVeSDllUodnRCBosEloDIx6Cc2k0w3OHBEU4/d9e6
Fpk/GHJaElujHQ08pZ4zDAl+g0mlMECbqoKqhj28PRpMTnK5T8eWGxm15aiTZdSLCOjE6TKBuuOf
f0KYFqlfnqM+LahkarZFtyTCNDHm3fQglnfiTlI1lA3YPispHZDLiGvQbUnRYycQgX1qFP+hlJ6m
gd71hM7lVaUB3K53VfiRvIZEke3EwKQZO4gNJTMpwG0zO/GyJkKjqCi1LlHKXWk30snD8WB3mJsI
qwtANTYz5c4/5VJRJQwuy6B+1WQNbQTo/T1LDskA02s4N8zKafojlJ7zIYKNWs1O7mB2a22Mkfhz
uJ8KwEJhmDnikpJQTtblmfIA7KW5D2eyqdS8MPanqiL2kfxr25cQtbwKjfkm85C2i/8gemMU8jK3
gFTejoxoRqhXmPrSN57qmwoNge+l0xeh6yTisQ86NV1I52w43GIYw8cpyw7eQS1j3jVv5aYJzF5+
aeo5dihM5NwgYjVDdOX4ebVIhWPZpo+YdcN0S0sHWExRik/PVDeMdIX1DU4vDHU9OBxPI3EFGFtA
uppUDz+tHdJdNHWP6bvXoajPWaxLpJIUCJBy0lrZUQS2KupUNeDwNwsrjhoBoCUGxOstjdxvZKWz
guI07ZuoAFHNTXhKIzROPfIbp/GYIlBXIWCCO8MNC1fFCHezRwr2FSS9A0+xROtdtIXzTiPtXiLQ
a2NVv6LEbmJ9C2GZpanp7dVKemaOlvE6czf5WROc72rfHsyg022PlgaGwlzQ7KFuflj2Mne8eAOP
OYV+6KpmAZiegC6o7XJ1R4AZFRX0yvtirgtJM64Pd8ph+7LSdJl35Uk6Tcem60Uc+hLYv0HsO4Wy
DPc7nJtmUzAafJZNiYDMFLVZJ6/CqK4DKLukcAVDu/KaqAibVjKL0qZ5045AhrQdg5x1a8EuS29v
DQSW4g6PZH3SNuZopySD0Ig52AnzM/LiUUWtnG19mD2apr28V2UmNsMDMjLCQlhbUSk8kCxNKbJC
ugdofF8ff76/gHpjMbkKrcRR3Zxx3S5sUGnjfaO0G8R4iJyYWIeyv0+fLD/6aru3cnyssif9fiNm
OJ5v8LCJsAbcEb9UnIdl6T6bOlHmKN0drPqt93RvZMj6R2OGldD4wqwbOOrogyzqVLNt8kdl2acS
UjSKKT5haUGRAAm9gtDDSZ5thgScYXGY3bpNrMBDOnYah/OSxdl8+1LYqD6WzZJMOvjJbvJ5F2jD
TbfYmfoNknm6Yc63tq3UwgZ9I4tqIgBAMQ1IsH2GaMB6QBj2mDTc2Gr7DgZ85pSh2YvyFe80bQnq
lqlrtuGZT2MD/yqg/2dVIKTBXhycuE7YRxmgBP56htBAPq6Wy4oWAYSIDLX+HtDdvRDSe68fj77o
bAr9z4GlFz4OJme+WcNw/WHko+mIR0e6cZiYqDiY0Fr8aOKRgHKmvHIB18gHMtwWkqBKFZlzn5BJ
Es/n/IF8Nb9IgSak5kCZ+WnQO0VjfNTMJZ8QsHiCJJSp9ROZnFFLqKYxs90vq83chCwgqQQ+FXxa
Q3GY/OjBQOpy1PK26QecENsZUv/tltSeQs7+U1tr6+Io4S5mJPnYck7q9MoNcaunA1MTRazXRVvH
MUaAZLB0HmYgWvjteBcpdd8iAjJI63CJZb/C1JQ1uJCdNOKZmSiHERrfRQT4UlARjmYMxAUnV8DI
jGyyD7lyjHiZCif/2Z3gTPyLFybC+qYPZTtVzQvlQez+fcOgoKRomncIjLkkgdkPZ4tudxsgtnU2
Mj/LXw3h/i0Trdm/Gqft68l34fygies0Wpi4gQ6VK/tXjB2xFbM6J1vj+kxJcdKBN/tDqxbvRizg
wvhB4Y9ytsvWMlB0t+ZTpJsNlHUpG7jSmlXgNmL6UpTCw7OZCOoHrXvEzczAQdoU4iP8LlToMSUo
XLoobj+eqM4qEYeZihBaRFPMI4ifUPZHM89f5bGUkjvcXyCoCYFgnU25j/Y3+eIWe1txksevhuRV
eewiiwSatqB8/psfg32LkcM0JGaZKSj8Wk9IAz1Hn3Ct/+ZGu24/UAub8vCtcFhbmtZihWrMct7t
Lz1fYaxnfVpkHjfkC/p5tCWr7ZBbNLB1z8E9C6ZARfl0uMvAOAqDcGzWUBbav6E4YWsjW3vw/Wfv
0AIXIFNOshGG2MMRjcsWkZOdb6MmL/aFL1EHpixFuu7wXCNsBQddS0UBy+b8U3p/PtgDjmfXNIVV
+gcki7evCkfsWMhXwE1tYdcAUW09SYFRCrR3isjMadhyJfctzBuXx/GbZOqjCOc7u8LtfwR5IfHM
z+kxCr4+/3aMU37miivmGYU/OGF/Ps0Bv1yRVJfG2+AnKsng+Y7R/5SEOsTTEVN2hN3OmptkCzrD
X6OupNT/UXFYBC7Z9MJzNs1YyQ+y9/x+AA0pQykRFyyJSPYLSQZz3Jzl5/rnhDrn3ESkxht47ecF
caASWsyyp4s9xgXJMmaBk59RrpsCpgAf4a9rfznNRn21Mil7vvBpdllZu1DOTlNHucuaLemNZT3V
VLYbZIgXjhCeS19PJpGwRPOYDTcy031z+zqosa/OGmCbjm3knZ6gAzRZgMtgRtys1DXil/ty5hkd
+wpGKyZg4ZCnU1wV6iDtEKd3b2gusa1osTjn1cHLIP8unxXxzdBpwsdVf9vRFaC44NGxF09dh33J
EuKj3tyHCw9o7pQV8TKhxyBpCBiH6nmeQ+gKQZRDD0zl5SwUk4Ip0DauGkmS/z0IOAFAZZBZnb3G
0RpgB7KNsrsU5Rgen1EFfbWTmxQGHdUCLKUgNPl0mPEIdrcepWfAHIjPyALi61mWcJVzGcKbRLRh
3neVsgHckk4Ow1glSMl+mfxBpM6b/OovqluYofSZLNQmdnHRYJGl3BPdXpCaKCGqGNtrG8jCmruV
YDhAi0ZTYn5DBj5bXC0gz2dgugEGyDx2upz3mLRj3+5FKvjqsnf0vzT5n+DLDBARow0ZZxChY0sT
SiFz7ISE/nJDxXcM/cl60uWhqg9CHfc+noEzFh7LdPa9Ys+Ez3NufIsx8q5NsiV7wARAN3QTTe3a
8f3buey64vJIpiloJ5CC0fnjLY9fOhBRLhzgTuqqPBU656mNOfF4Ljq+OX8ttZ0lBx7k/BS7nfW6
7eeWFXfZZ34HUQ5iWcEecmgqGoDLsR5DBOc61dmJYD8al9UZ8cyaodX0s+8lM3Jdk0GKXun3CZ0Q
7TOhxQ3vbtg6eqDCgt2ii9GaLEXa9+9ciuu1igG7yPf2wFtofSLtfqqAi4i5S+mScu/CaOTMpRrD
opaN+at0c3IIZ3Mcu1N2j6srd6+64X37FewOqzZkC8nc5ElqKPfSzbV64CFgWNyUdpIzFVXoUoRT
iHY9xbLj87lu/Uk9DHRO/n6Rq80Snyy+UBC7/g+I7/61Uiu0McViD2UrzJeCEIAfEdzcKvr/behE
zhxnpzuPCxOmsuoaw6w84kdV93tU/SlcNSJQYDlSHSlFUi2u0QGj8gCGfnVXjxesgDJt5+mvOcfb
jUaBUOOKIRsxTQ0lf2sCYLKgWa2+CG0OacK66rZWtpMwYqaUXTtn4/nctmV87b8x5RiBZfsrK0bf
JChnNSQPHYB5Q2wBS5blWti6z+WTG9ZDvG1bFZxh+lcgZYuOjoJDAkNGc87qsRI5psgd26JOehZm
xC5gfLaRc6/VPLopvUaIO69F38OyAu5evENcAPgS22kxrhNzTm9rT8paKyX2o3vSzNAiW8mO22Zl
xFpHv8/WjyGgV2VuhvanOefxTkO8mn3jMslvCeau86Kpk+YuGK9hXrKwPk8QI1Fy18g6gJTt2g6f
r0jJvRUuH/20MKVhIPWLh82gACxutRp9xmcGtAJ38X2UsJkAR/NMO/w+VQL45DijUxQqiJRzXljM
r8lroDBV8Wm+H0s0q006K0ygNUdjeizTDgaXEsP9PGO8oLM2pI/RIBlTxeGfh+ocRTuTFyaASJGh
UFsboxEBbzvTIFxQSicBrV+a+1jkqWa4NtuONM5pLzpdDodd1xch7H/7jgtmXQiaiDf984pEERRm
mxCXmEkjfD/JUAZaSWyw4dw/OkCq6ETuWQYh+axvc8Q9o9zDiyHK8UejfeV9WFKIyzWiRe6NydjM
ltwGtYD8/CYdx0vMuxvbTrI8LxMYxhb6DxZTeyUmiG6lZdxqi5qq3odfZHOlL6eGhNPJ5NI0DXom
ypmBthvQ+hQEpBJ5AnShvNWlFtpnzM9+l71jSmeedQw8kXnoHBsV3DqQ4A2bWdi7aN/30uKSlTeg
VfJ+qQFHIF3hUfLJl77bc3iXetS+BUzeVsD2mtPWcLcNYrvKOTpvlc1chyR9hv1jh9/NpRDTpyBF
clOaFpQCy5QxLbVJM7k/H9D1diFOiBLbHDOwXvachDq3mggRcM1iOsEbUzLgxeRS2PiL5HC7Z6cv
TLZUMRtGqU/9SxMQhc8pCMqbkErQTYzr/0QY3xiCKOByyZ9u13Cy/OJv6JwDALhNdIDRy/zESoJV
nlDY2l4lkroAdsB8Xz5/djLOUVa/v5QUtt9ewSNg4TYlJDFLkFP46b/T1mKL+Q/XRhjlb2QCZ5mI
IBgitKShPxjYVDNiJuSWt+69IBtKCuWoDTA352tgiU24twoMwNESBfzDi+AtI91aisiSt6ce8f46
clkSkVzck5vHwMcYgHIU+xYlAsU6ICchNoB33QLCtLSxvVkQSw75Bf34iTvSzgqkuRKUF6+qnE/B
JIzBMlGiLKt5/2KDrrILpQj/z3TfMFKRz0jdpbn4dnl4L5UE5gY4RgKz/dNSVdNjY5LzqBliGPuP
tYDGnHzM2718N+i3f7a9ysrxIgF2AljO/++o9R4MKSqh4YbbA40cAkVvYPeji7lZvL8Z3cZrkXUA
3KPCwJ8ZHqcGXC1c+k/7fdJH4FPYSjRe4+YwGh+acyDWkn3qijjUx3sxEWC2xTBA1O8cxD4elTa6
qhMfPtDALIobWZxeevSnJr39QOdsEZeS3k9a+t2oX6oeNA7Ih32L4Eif7J3wskLoOGy+xiwm4oZv
UPx67Un0jYEU5b8ky7FaBvZXwHCXhK1fOJ2NBtnzGUeahkqMmrDNFW9deP03Stq+R76L0rUR7DIH
V8LnBhloan7Ut3zZK2rNCFBTpASsbc28kk10Pn23se2ZBfABFOJFgC8Qyhc/Zu9ZK0CtenMJ2nxz
NAZkcbx4MKRYjkSnDMgge4r2SHYu/XeuC7jE3L85O3Jx5v14QyGjCO5+UIsKSlyosfxy0gJyYgVV
gkiMVSzU9igbtOkvXwMn4UxLpdnGjQhBsOWag0HP3Ey8xhagK7BdRoWZHAFsTmLH5uwQST5tUvyk
wiSOtBsbFw96ByUdIVT/dPwoCAWP+iXFDEdjAdma6Xd1GuJBTyU8r9M+StoYPeJHTgIGG28GzFQ7
Unpr0AK+WiwOFVSlsm8i7spKSog5BcAsjt7yyUmVSG8SfQ56BtXZIKw2Nf+z7+5NadNmOuKC1nHW
hEifYgOq0hPuKlYWaMyHldk21rxu6QsRz6XfGb3kHiibBx8kkk3Cr9JPrGAHhJGvEbnEETCDmSeS
Mlv67KpUPL0Dgwfhu5d948s+N/c+QVuh5oe7KmOtx02URjAvX4Fqjn/IWJEq4hqdc8wWQrFmWJl8
yFNGEhA6rJrIUDOxT+V4URmpvwQHP7vT9f3Xn3Z3qO8WAArhjt320Rc55qP+5GgFfVmVykf+z0Eb
9DizLFyVkQ5LChx5ahzBCQmccE+fUeg76tNfnYBaIP8iVHoXFhVtWkAiOL0LwEX9BpxNQsmXs3S0
BSJHuj4Wgtsc6NmOhiTpEvTHZ/5YzrPp23QkEJAOF/vg04vOTnGAt6VgufPoZnf60FB5lSFazhbd
rsJmUIHOlIYJmmTPamox9NXEFJqShb4u/LxRaxDJEr+iKxqyUoh/yekAMisMF604ZMdvxxB9vFT9
koWXFa4Ocu6Ey0JhCP+mJEckeBv7uxnFFoc78RM4bqHT5tNba31ML5xxRq6FYs1AkxEH1C2vAMdn
yvm+DMhxUta/xhUuWT6oFj02da0ukvspy3hMygaqJK+b+tkh4A3/akl+IJpOoUAYJQw9kDALqW3j
eykZVQZy7JOa10Ck1BDhWwUkRP71h6whkK5tOgH069OW/GQ1/FMNk8vBqklJSKrDRgot1dwpU1HL
xYYl82voJYg1HZIWcYdbaqF46LWFe57HxBa4arIjKvOemQqxl3JJH8VJN3CNrSCrR58Dqrv8iVUE
m1oexKH4BIQ1U8PoekZCH82TVApM5X4yNxDr9QkaW8b4ZJ+zRxEWZMgkqWOCNZCYcrhAwsTbvvgg
XDhb0KHsWhoV/B+SDnnGGKyBW6LQhy5hwV29ygSppCRwQOoON+zITec59n2+oGd6uq6nwh5AOC6c
fJDcjEiC33qxCY1Jn1lZ8pUt9aEkcp6k4DGxI1Pu16KmqVfRaqZM5/JFwK60cDpNfcTVup/+CS/X
grOz8LTo8USS1viIDBdGY/H0gueGlh64Qm0gVgCu8+hNoRjpaAU2TKocUU53HVDaUTN5Kzq+SZuS
bk8ftIDePRbEumKS3lOp/YkNyh/hYlCCYBfi2ikcU9eDJgalRGn18JItJu02HlaAdi6KvxM1S8iu
8hqdeddzZba+Y33lL+xEvbngaTpSi0N7Xj851kSWcwcLtNE7FjzLVUpdCLFpsuX93sij8p/WsahQ
Z184Pexg9px7UyI/qrHBQyIcWHRTGVbBVikPJ5l3MXcCaeA1a3YT2RbjmdTz7G6ADdBWuXUGSCOO
p92a+/4NYceLegsrbjsweFkJ9t7x1AFkCSHv/AY5FK6xEpRUTiwhIv69ObjoWXEfpEdQNLrB+/CT
1lt3/fhgLLvD5xlRi2Jk3MLTe7sQWTaHvU7y12ecewiAYYgrGosKHQ6spDWaJde7pqNMvsoRqZhC
nCBbt5MF1C0GQVc+hQXm08FfXhoN40BzJpxVt8LL/WBGvJOzESvbmYBIq0+sdPE9wWJ+C2FaUH+B
fp2UZcOqB9Mx32AlydWfl3Fs+EMYjP5PgiIUyiY7urGh5p8iOj61Ul7nLVbGI+kUGKzM69ppZcm5
0nziDUkaZ++YsroHVQkCHwpT5UAhmu1IFYBFTURGzbzMpC0CMu/C8ji0re6BxUalvQUnAnovMPWr
+nF9MBATf0mnrw6UGqO5GXEx2e+1rqLdu09jVK9UUn4hm8lhlijFscnyqfx4lE0xn7mPkBg1awAA
2XVHVfEMs0szakeno7vn+wvHDYstT6dLRwd6PvkK6oysIZ9Fz0oMNqR5D9b0VHhlnhCmcQk54w11
LwCd2aef9K7qZcAacj8z9sr+wbRfCGdSPo+p4ACNambi92pMTKRI3yAEIVDCYdL3fgL+5eMsiIZm
c70lvdFWftnw2qHRdXNZB4SflnQHeUZRujMT4uNn6HQcIXK466GCrG0uCRQwilBGiB0qE2mJFMxb
o2Xt2UxdUqhRE2acUc/BM9F0pYen7w3Rv6WtTK4pQ/sA/fKPzIaJOqSEWzzHe92R5JdTTfISRPhr
xIyNHTwULyB2EIhAQxFd0qkT+v6wU63IFzkWse2Kkjw/1C+crCaRsw+/YAR+6ZLB2RgpGNwaPaQk
cQQPuC/O3TX2VBkZqheNtk2ZOdWBFvJozpld5UIkoynLQw+t5cIK16DUcoXnrLIp7Wqav7NTWL9q
Yd9NsxTuFujRff8EmPY4GmdoSe1Ue0zLFrf6e0i7iSuljr2KjoZe8q7GpRT/Rqd6Xsmqvaow/8ko
AA09uT1mSlrrZnVjhG9dnubp7+tlVQnzKQggZGDZfN240Q0gJAs4nAMPEQYJFUHKSlaeQKNzEJ4T
CJwfhTHXXbNbjSzpvk82CN1KT72s1JVpQ6jesBA8C07I3V3r3gOS6OUecZhsqYi/Rs2GkzWJy5aO
KSUsMx0QVEqzoyuH7TwTDQTsdi29J9I+3bFmadWxecW9Stx9D1qju9YS3sufmKTddfbgsSTOk/+M
/QklDChBnZBF9K8PqkA9OW89ZlRvzlDIZfUbtyYGWaJcm9R3+s22lqNtrgA+pMS1i10W4MRDwRGH
+t0KEP4weFIk9cpN5OYVSbY5VhxUArpjWubTS+PzbGHDipy3IURtzkOKoM5hC8RIrGGDfJsDd7FJ
fqmdGfGvB+HOvnLWyxBM7eBTGxKRY3py6M9SplbubQbqOc0GNTFjmV1RlZBP2BdJ/irLQDpGMlYg
ULc1OxvgbIdljHZTg6YWJ4RN721Rlz5XkB9KhHwnI89DmJDA+9LBr2VviZ1izEWKhuMrZxnIYR7J
9TkDjp8aoSO+G/sq1BT3ZgYl6lWbPMbFusG0pxp0tvL4mGlfFjA7VhFxXqaS2hbBWHOEpbJB1oMh
oOIUCacGRM7OgCrKhP4One1CJYOcwcl3g6nvg9CzDlnhpyVh9taar9NC7nlBYxUDRtg+bTbTWWJ5
opgVqdSKwQJswUxhw8s3PpcHcv3+29HFo6CKeqdW4secncQteDKqgc/0B5/cAz8DJQsnnA1zASnt
Ekb9NuvVDwFLXQJjOGrwjp0ThKQsUOUJYm8cn3o4gD6PmVYgVq9v7TgVr+3BEXf6wsrleBqYrjcO
5rKpZqTiF1Y1VTYjXv4vnfCmgap7AOE2q7j9pVdcob81+DkVR+8LR1Z+5up0iEtptdyKauMO/I29
9ouFBKM8Jg6Hpj2BHlo/Qblx8cc+hgrXVIQcM84ae3vcpunbceEUWgFope4W4SBBMRH+j+ekR+9q
F/JnrJw8Rx8kkwI+QEcLONcUYwZXsVjYfGSm0rT1r/FMMyCgbZEpcPtRx3T8hVygXqUVWsWc1lWR
ezLHwb8Oy4bytI7guh2+PTo4RIosDmVzf+r2B3FZy1Kn+gX2IfnjPIUaAx3L7lY9dbeLXcoMq+3c
Fr49XY1hwxE8SBs0umeqXg0vToBu/pUOQfEvW6HGpN+day1YiFUH794XmlD2yO+//6nw1Dvx1HFc
HICd11kZv8yQyRZFnpE2Q8zkxImqNVLE2QJqPQ25/96BEjzDaAjWbMB68145HOm4VIOY2bBzAD//
8CJ1mDbz5dVJkUcrX/9Nly0usAFgyyEYHblxwUPfX2m95lVVVAYCAKlLUVVykkgPvhlzqLHXAh1j
dbCTuwmBD5esW/MNCSMF+WuhVDMZN3Qr7baMuYVaWs8OiNcYqhdrGRjxQbKx3O5rTVwiCWC+jALe
32TziE26LGF+S2V0B/ldK/PQvznNEy4Ur8BVD7oD/8B0PaO2RTEc7rAEW/Y+tZjQGo0VyP95xy1A
8FW8wVounBMywwL2zatKFRCGvwVtxSFHIUCVacJiePENI43k5M2skhWnMDs29+ke2DkuZOw4RZga
g7z0vISpS3fT7+RwiAHoVDREJsoBUmnO56h2jExXuLtxovwnvIyR67JDe3P6/5hAqLp0kScGSfKS
zLHKiumws4o1hAyTJnt13aoenapmT5/dRJYa3HlZEg9YQ1hZXPrgSgM8E7DzsWr9OQ3HT7TBR2z8
JwBjJK+bLKwwnbz9f1+u2CR7ucXe8sJW8Q3bPtP/fFk5IFhA+lkozqepb2XrGszVfFzxFVxSJgAQ
Zw9SpuLURHGAPv2lJEkpJOUu7d4Z4suliQUgpNSCL+SPph2oB8kvp+f5ypPjIhoFP61M8nkZXTbQ
YtoZPJBaEZeUVvtEidqhmfokfnygVY27PZtduVYKUtofr556H9ClLyrTJ1kQNN7VA8KovroK3tdb
DXDufZArz3xhTQkaYlRgvbo3hSVfFz2sF8Kxw1excZqUkuehz6iiRMBYyFRCQ6nRsEwvKZWUKuNv
I7Y0R9twsBQJlrQ2r0AyACtRERkFTMpk5M+qSCYTCTVELP6IXBrtDmRNPRuavCweu9oWXdXwfNjK
sD1kK6+hv31qp5XBrDCmBkuP8raMsr2zJ1NhISj96u0z/GrDthC+592I4E7G9hz51M+FaDfoWWJV
Jtv1jLBQZJgLFIC1w7kB/MBWRJ1bfCbr67zXv+phiwTxNUKeLGNzughY3lnQKk0Sf1dI1zKwEbkx
6bCQjji9EN6faJw+skgAmerkDMlYj82aoMt0uv72N6u9CPza1GSGJH8+aXsA104EKIAb/6ZhXqJQ
BbjPoIvaOUmT7fyrW19Hrq9FPxx0MDGMTpyAYGgx5HraGAQ5CCfSdm8ibNuCwOo8S3zFUhV/uQFD
782XigMAHe34nD8L9vv6cxHBDXsaxVEZHrdTjl4uQL5q8JmLYBwYfgVIg7rzrFqJZStMhU9aDyOG
3il8o4sjJDYQiHHKeGgnUMYzHQnwwIklYIlY6zExd5n0jjtUcHRBaH73CjN8bdJINzNabZN4zScQ
W6klx6B7ftfSEmE9YdkPbUJuJSZG2wD99kcSKI9+z9I5cqNYfObGMcnrQxVUjpiFrPJnTVkCgzvs
zA0ZsNURdtO81iqHfvApvne3Iu4GJiXpnxx7QaVZDPGLLohUZ2VFwAsi8l3P+XA/1dnRvf7zzCPg
tsKogal+chczfJdCglg5CTij/zNv5S0euqRgV88fYr40a9WqLxZQHs9NyMk+qJNPeHlKhZkbQqBR
VkLo51a6nAoD987GHTIDNd4DRuRiFO7+13/cC7RIKNMNCJ74s/Xyv7PXn6wmW+NfghXtaGR6RRb+
ckWO7OfE264QgljxB5GdFagw6m8FB6b3B4ol/LtKE1HDN9aKnRpyy8BDPiWuHaEqvwoH2Ey9zu28
x3yIO41sRcaRUeKVLghG3Kf0yzVuBd9weJygU/tuF/Ogi0rXcYYi2hVm7+CwbW9rL1uv4bPxATOO
xBrpBa8JaKreuwfvabc0VcKAdW5KxLDtg4gAAjcDYADb3PBogJXSssAXiw+jBIKphP2m2YtOaUda
4zn4N9gZ/y5VFuLj3glHJyv0NzNRIF4dfZ0alVDfNLpWEZRG8McyNt50ZDIAuEshGGLVGa6KPy//
d29998OJPB/RFNqPULzgkk2iyBEjmww84QjhzLp24lHsy4uoHZQnWwFeUQQOMi+677TY/cqIs9Cf
04afIzDkli29viplcFTMsQJ1AIb6GZZv0z6LPN7IkF5xsPLEDY+ck66kPXzJu0DnyXfdZwavZ5YT
N5X1flrFGG6ayUCaURqoqdXYUHQeTa7m32YjxHvsCWzzYh1H0b6FfhVTnCvP6BMydCX4x4PnxE5C
exQgghMavFWljvDTWahfzTeDqSzz6esqKFeUnZI8GkxwiWuPPwxHzpnh9rylaRI5qV+Q3k7OuTi1
8+t0fKJ9JMTSK9buaRbRViPcKkI+o5ezNol6qS2IcvbR8tWPdS7LnAY+8WiB544o6UVkB+DWwXa9
dShi4OZnOgLEUswlH10zQdvrB95P8JfbwZrOtnLP8IaAt8d9NaptVk7SKu+T6wV3JRVcMWIs4mMv
i3zTFANX1m4/2EGxbb58+fcMu9NX2vU1Xa5Hh67saS/A73gDh8d1JC4f73zatf5/Fxndv94ubxKA
iGU0EGLXuVRooGpTfnkKuzS2IAiDOLCi1H7oex2FZNoJ/EmULEIGgRmd5clH5AZdzLro9XHLFZDW
W6t3r/E+obzPErMr4+NgV8flmFOt+0mcueWJg50+b+Nkj/7khHzO3KpuseKk75TTi0X4Ehn3kCxa
lLYWKPWJHFycZbHKxqJEvTVKDWd7plGgeXLoeGSxEQk/8M4L8tzoYdUorX4vqR9RhwuQcV5gD0d4
zQgSjKgv3qBnBeca7/weYxooVxhbAuAm0TAV5qUrTXP90ntrQH/PJrpI/Xkh50yNZW+IgtVPTXh3
h37kXUGeG6LEcU8HjcWzJQ9H5DS5iDsDiMPgYyO+iyLgA1zg6Or1ElnuZsJKagAnDotCOkDuA6ip
HmUqu1RKISG1Tc7zcQ12Q34XSVUrNsrMov9JxJG7baCzwdlW2WzTh0BLF043vaUjZXcpHQ959mh0
USkZuaQtv9lQknyCZD7QW2++99dJSPAKGs2lIMMXgomfiCXCdtEqZrswBNxDj0xdhR9TH08gBSK3
gjdUkUsG8298qr/31yrkOd7nv41sSq10GFFfcgyXTx6Mrw1wzR8Wh4G40qw0Ge95B7gcsrX4bW7W
SZJpfIzP3eDM86OhAdFjGsXO5IqHHK/S05hnOmohPPT4nV+k7NYmrgXRtmnQUdlVHRjy3lzc+CmM
8YTkWxceV5iNgCsp/fLO50Ik6XOo34woeym+S+LbxSKUx+xVE22Vzm2pP/4zp+KXr2Ej/7KAVnvq
V9DnS7MmCEWR5ctt4Qa3/a8SAEribL+SRwFXJ+U7myWeBPesFKWcXICI04WcgWejUX9ijBQdQ/qj
rov4O0F0xOEIQVATxVkywTcS+c8OlPqwVEY934KzGtIr82ld3GnL5AkY2C4NqA1oUZZWPFLBDGP9
w6qboqoj14MkAVVc6UiDHng2120/PGAm/gHQ2ou6zxYGnMchuq2TSIu5xivclzOFnYirUHQsJm+c
fS1D6TOm3hc5pWf/OBhyVZmKYo035I8kW4JCzrveDhxxbSopamdmSp7TnGhCtysVbg4q9W7MXVbI
l1TP32r/JFBFEGli18vgiGqJyMT+rgH30VaiNC3t2n6gIB/louGZ4Rlm2UpSHsDFnwSHG1igMGh1
5SUJrMiSKUOVkv0+3oUSJjUKsTuPPn6Nmn95wceoPVuPkWSe0tATlRZgjjZN7qlArYt1cFI2tdUj
zzjpaoi2qi+XmfBnkYbhTSJ7RHDO55IUVIkZs/zX4WDm2qzDkevzhPSMlckbpJ7wl4k+KvQnodID
M/AfEU2oz7dWEYm0ywENMf3lPdzTyoIWEQ+OTgxlvM14MNmoZao9YjMk2X/dAXOejF+rzu36Scgs
6TBu88vKp6PZlsew0+/VxeuZQfp7LGwKLpJ/rsCOXS1nEQ+bhuUY5pNyQ3vpXgyoU4C5x9BLN8vZ
6C4UygcKjQdSsgIVo6a4Mha02MszJAveDIFVkR/FxeWPaKxlqX02XubgaoyqVifMIwvYECZ+7H6L
KORr+xZb21JmKc2v1Sfn8aJl88d7/BxM0jtd0oRtd9Q6tzbKbg6vy049XR3KkJykRgCjmVRbCLbg
EhsTJpprcIlhjo0IJw1NcJUsb1mHL4PHy8wU0CPzz3qtCiCkMs00pzUQNl+93+7LuuCbX/DGL7Px
CAlALff1vhgZhBv3klgPzi2yN6L9O7ktOKKRsZpcaBaaMos5N30L3theoi0fzbAtc99FDHISlqhX
Wwn0CgGkACwqPmqcDdvdIniYn71nnlQvbMBxnrako64ZF/B9t1DgmV3i7rnhQ4oNzpZSsHTJYjC9
p8fEQQuPrIhjPfjbrBsAS+jBqfmWqRXjWIs4cdyfGjJJGFWGD5cnaWTFdmaO5YnzzQ2rBIhH2IBV
Aq4j0Fpvwh4OMsHArSegB1oFw26rGYFvA4gZB2H6t0lEx+A0Ok2ZYR6UHG0Y6k2l4nUPFru8W4SD
RZFvGr1F7Fi0hYg5zUY3Jb+RCPDHeDtbRwwXS3Mjd8PeDDBzuC3JPkvFp1v0kk3W/eIu0fn4QypX
8WESYt5/q4CI39sSHlwu7U0XF0wMGVEKj/p7+fKjecNYrzfAHbTNrjVyLVEjYGx5Yk9YjmSIZrww
1JE1t2HmscsqS3lmdKChyDO70FoxSWuPtuYWhDCZJVGD3DVvGzKL3nLHef/mElZN6FW3JNuin6/z
4ZIfVhITexvw8DVBWNvkD6ZmP9O250Jx9PJv6iYj6lRO0+/hkhAUXmc+r5NzuJMqxzMAXmhzZwsl
mPbqi9a/TcJE0VTHZvUg7zxaUSN2lt4aBEcSeVKDT5ZHs7+6lfPvGINVkB9T+HehQ5emMAW8tnTy
5V4lQ5vfy3Q7f2MIr/PdRCjshtQMY63YAyo9/1PVhi1zXvQgsjUueXYz9tHQ2x3knih6CL5SD33n
mSLDRMZZVq53Vxxmk3O99t7HSEMkMRsHWxPh35hM0mbsfhuT0i1UIhE1w9798CGA8oQgDd5A1ZtH
uOjou1a7dQvpN7lCsCUCaZMRT5aISSZfm3I/5ahD/AGfvm+HiR1MbZtaMi6zYBdyX93Zhdj534FB
MMFI8S2HJJ6B/mxRnWLqctFtNcl6GbO7ZRnxKGQIvWdu6KXuV5MZhlMM4pVO+58dgZSNNH3PGTFh
tGOj3WSPwmNj5z+A28N5FP1EltI41BbC3sKkj+Jyp4NPDheotLr54eJUEN9MmF7rQtX1YDntSwc6
LZeRc1uyxopvW7TwZbekhf0z6a8lvZMxT+u6ul/Mo/+YiNHRt5yv8LyNVNGXvd2G7YPHt3OJ6xl5
t+qIsycE0cQGuMqq+W6dxhLkisAngeLbxY9AnfxwQ2pJOocOGgnROtcEw0UKoLD+h9gml84Kg1JQ
BYHrQFf5fdghPrZto9vk/y52z22153Q1AlYYKGXA1lG2+nUL1N60VFweoCbQTXFU9w2nejsM8QqE
LwKmqFrThUaY41yj8EalwIcmiSedQobVJRg398fp9AA8wQM959NC5PVAnzTvpupTZ7gO/lpwD7UD
tGnoWd1rEmBE5PM9fq/dgHsxmcWxjCgRe4Yhs1H+RornUO1+A+fpQnegN6EQlUY/bAEUr389Xsj6
1DkjlE3XGGXhFEaMB0/m4z4sZf2/zeyhSuIG0hm8e2DMQCStRnJpYS1SmZwFEGIN1DQjkvoEiURN
n3M9nRjyyFCjypJNIJfUwRjy9joohg0Ke2om6iUpFWZC9bJ451dGIZ6TSps5ziIOLrxDfIAHCOuV
A7NAePx473FEamaJvFHjdjwlkeuxsXaQoCbM/hBR+afCc1bEH+45EfuUNo67uF6PgK5g1F9Fy5un
Yu3A7fW5zSNnLlvuBs4GrYOejxLkdLqPttDosPkH1co780XagAgAM+JfScbJqnlJ2tHT6qT2Bhsi
7jcvxmdX/eskuUMTUI9EinRirt6KukYnlsuK6j/WJgzyplQOwWaGzR8lEUHf2NfN2s/mFx8VvsrV
MBiyg3181FcfGSHNZdmcUY95LhHu4g+Ajsr21jn6xyhUf0nKG7+6w29dgk5pQn+yVWTD++kPrpT6
pKrUbA6kIiMvd5hw2u2ySGh2yHQqwSB/KJ5QOnyT4egx37Xk8lkO25Tp28stLcUk+UFnNPPbPSg3
jFkzrceJs8NZ8u4l3NCt1D8ynxB2FRNvGEDZ9UiLKGxnS3acZFLKM5DjXp1GIvFAD4KELtJi+c23
NxZWuk549fCIdEfN+WZbHFnqLUcMNozgkpJRuUPPw2XKKsB+WRJbEyq96HVeuY/q8uFmDacGFcNC
M36zDuwn5KXbQ2tRQxyZPm87JjF0uWqcCefugoudc7VfAYNWrz++vp+X9Eo5uTNfTOfi/x/s4kIo
NRJupj+uDc9jbBl9O58Tk+rEK/iiXh9oDv3MhWMQszd/zim0b0zYd5hlcKp/IohjEkmjXa08tBRW
BEZPj9c1FkBpecimU0odk4tU68ueEFz3bqUzOiQrDEdbTjIEHf8IQx7AVrfOG3rXBWTiqfL8tp76
5IVOLPnCUEbPmrP1sGFx90pp1MffGaQqqZRa0CJhtaFx7JT4zdO7OyWds/U/VunPkJG6iwsSQq80
hYT9r86lDA8exQsyMuixy6R3l/HK4Uimwa+rLm/jW1TgaTf+83eT+A6kwV05r4QRkDePr+vvIoq2
HM2d+IgowgyZj9Y1ZlYochSL+PK6qK6F7ip8HfzW9oyyiYNHQYuFA/GxeMaAUaWn418Qn6811GJm
CMc76ECOeRtEAlNZoNHOBLn6qWCqaYtG3Iy0/FtaZgcT4BIc+T5JtN6wxEMTNVFWmeDHhx3pHgo9
zycb3nFAUkcYkN7bElF/aOV7yvWFlkVScwaYrE+HudddhXfwRV5ofan9TCUOYmohyiZzC3FCLQDm
TtmJVQMc/9irtcb+0/4j1MSVIqd39RkbJMjFZZreYO3L2/ZI7qauDpeQx6yF4rASa2K3IS01zS5j
hlCmHgA2uXnPm8uLJMBcoYI/99uozzIvdmh/oXGeaxQON8UEyY8NNtXbfxVsIeOXZcw3mRpY64CA
Da3hsfVhU+2HlE14CDwLDJM1MVjtAeXmDs6TQeq8GV4bczcO1ZpOq7H7kzMW4x9Jxr8+i1ztMsui
FW+Wf46wkpQ1ZMdqKMqoBZUg3/XPqzoFZfxgTlYVNAol2une3jH4YulYKgvmf1l5jKy16+mJ3VNM
ddYWzh0J3tqYFzjs3YIA/t/Df35KSviQFH7i5x4aTOEgAQ3gV5q8gh8IT5nmwxRubCj7HOz6490E
/OOKL8eWWwTHvWRTPXmgebfM2fIcTo+GknvwlVtkgjWKw18ztABPeqE8HqjZNZVKKmMVpIKkwnjC
g2Bz6IfkXJolXwuQYw5WdgUqUe8bH0/Joy6UMx8BTIYEIfE+KA7O5w8yTs2tQuZ+koRXmSo+Hs9k
xL7W3X3qs/GnXilNMPjo3Ma9z9iBCngHDTT3e+n7QVI9nxbq272+4TMZ9AOMe6Y7l8io0kTZ9LNt
7UG0ZtiTRtXlx/sQTmQFkXm21ycmxNnjDaSv+df54ZqnVyJ/ZbxanIB57dr70b8OzWWPkwXVgVFG
8vPOcyEIMTJVfluR1bpTd816+dyZ6JpBcpVhzeLY8CF2XGckc6lyfJd3yu9F8na1hDykos6Dk5ve
G4B/q+W87ZyrdZ2m05DSGhl8HmrLwfNIepqZTNpWu66cGETk2rplxaaJO0g65ekvX+IRbKXo8Ki1
UcQ4oflVrPZgzsdKdvwF6+hBSvZzARMRZS1Br21X+xP8/1UM5Huc7prF7+VWeqaGHP8ikNB3lDBu
51uxGNSB/6SKxAsNH5NCNHIFaNclzxDmnEQYS/xX3GySyHYYmYZCeOxo5/tnbc7OtstjTNJYg+PJ
mT4U4+QBdPD/PDOrpImS/rgPoCS+PNhTvh3mPPE4t6pYXwBOntJdZKFz3+pQyuIm+2/gUCowJYYb
dqLth7Br3VaTLijR5mZOK1lctaIemhAOZ/AOhYJnk3T159pqYDrZZNp4wUlwSPaRw2cKSQqPCF/B
RzndIOTcUxz5CRV5GtV5R5VS6fl/eAoiSsHAhfVancPsuuu0o406Vr6YsVaIB7fHDYfBj7ZxdIyb
QRvrM42ncy2NO6dESyZyaoocRgNsDm3Y+CINZnsEcVLO/vqyfGROj5UabFahGuo+lmy/qgUyLRY/
UNQktTu7cp4ttZ0+2eVL7RiHVEM0u9lP8JSoRsGYx+EXTYRvi1VNEqi951oGudv4fB6j8TtrCCi0
H2jPqhpJZhNwyLg56VH97dWplRtpJm5jzDiiUCoUfvAS8625jjbNcPshxfboX+frJSPqMAMNLfdb
oQMTPymgbelMlMnb32pbAIUEs0e1FEJHzciqHlL+FGwaj5H8fh9Zf9JhYLTYvjnqNqpAH9/ccMrB
rFDJv+7xqyar4gjlyQITaiAfmevxEHliGHKFzghagEAQIpG7IlHqp30b9HrwnxMy3ySVhMDP4Kza
tKzUttU9Hpzz+R7CrtVvAip4YmKZl8IB8XxSY28pbrwb6FjF3IOuOaGvENjSyqLKIof6/Ucwq9zq
OJHIObQK3vXL7vQiKeldwmxF9eI6XPLNTb/dJvFUjKbWRbXgcZ5mfrIdEBu/AgtCt7g5Jr5iQ639
DFQ4mS9pDirXxpDUOzlVnILzgQqHuAR9jdnHwj5w/acsavvdXa9rYZEkph2+ixZ5S2XNovh5QtM5
BNSfKtr5UPIggH6iOPKubHhrpci9LjjZ+hcxu45Bonda3XNYzFdTnfDN/pxonQ1SHDBkPbGlByro
btO4Mlj2Dha3jXigpGYtPtJbTVDpyeZLzk1iP+/wgvi02SEkj5WtRT/+AHDA6YM8lWOZ/u+MPUO9
riWPohc3mtBYLp5TIh+tULtmQB+QnNqA04t3lVY3mgx3P/zsy4waAIbUNAYFEf/iqDE9HPgCCjhn
HdaXDr/LaF6ZeRBsTzlLxAuD2Y3ECrfbjADs1DrYJvQ4/Icrh3tdtPW05fXOxJnh87MesvLWxtqe
Ek9c5NgEVFmtpDDfuJYaUKwt8Rrnts/YHh2ia1vloPtJGLO1lmLGjyvvWnnCvB5n1Hbb0sc/FyLn
YYV+3brXGpXgxNMK/1+TmHhAYdUG8+J+2L0PIfOmX5n5ZE0q30vrHAvf/g90ZBZWtHZESmRBkf8O
N0sIAVH6/aCTx8mwB1CMLQNO0CkY/aNKqxCWnOoeFcqX58ZmRe98cuQAmgV2kYhJksgTwz5zZ2d5
1mefDEAuuOYE66JFoURqvWmYZ0h26K10yXzZmMgvvgya7QF0sV4wOT3Qf24xkov9STVxirBzm7Zq
mSd9v95vTXvnkhZEIewxsIy9HSRQvLWOf44fSypLKYtBPoBsNEPfMuM7ZOf49Tm/TCjEhFeK2Z4O
Lut3Gw6hD1jx+KoZH1Y9ZeiVnmH7uNd3PG9oFPZu20TnMxP3mUB8HJfse1nj5qfC66m+5KkBLnxQ
/GdhObd4ZC8Hf5d+n2GTYmGpAZna0yvB/98L4SCyMttDSDQWY3yHz8rLvEWbal6kxMZ2jptWdP2G
bHCWvH0Fsp2UFZCHrb3BlPtP6E0IJHVGaVhb6suEEI++W+ucPcb4FbMShinNSxKo2hsCCFHcIeQs
bZTM4LyXu5QQRit5teYO/8e33KMAzFAX4o7EGXVTtFsFXpMYsHwn9wfITYTa58icWyWEG+3Idzzm
Cfln4dKWCZvAdOdeUzgeLbfarubenL4Fx4Iw2RgPov9nK8VMvD/7Fn4UxJtDKONv5ke6Lt6N8bCc
imVWaH7+nvQ50+552/y8WqxxCRkz7YFCsskd81hWr0pHD06aredd4ZFbWkyo2+49GwFfRspdlSLp
mAB0yD7U9zAdNp2I91E3K9DsgYEF7Tj5aUaFQrPlBRyMPrf3g10+bgMRzBfn2yz0OYFylkWCUa/P
ycxrhygkuK2smqeyfyWO3oxiLFjY8kcPjFoBRTFLTlhs16wrTGiv0/FoGV4OvPfL9MhQIRS3gP2V
WwnCqumV6HixHSjAVHptnzyLPH6xCdKYQMf34YGa4vYpHasEJktoxL/3q94rwgLNZpQb5Md0/MRi
vIiThiDHlntvhv24bzHWftdb1LMeSeGBgWImJNVfO2ny2RcB313fssFRYJ3F4TA78Vk72IxQavK/
I+qKK5eWjgcNYFNbmmKewdqF3TRNsjHDL99qvHCtzpswGeFmFUS8KcNtNLyeCeIGv5kykZo5Qmy/
puSLkFkkv4GKhOeTQC0Rf+3gkQMHdMqxM2lY5KAWjwQzP1lg+b6OPyyC7kcpBn6V2Ur4z2kHJTu0
uamXNmml96p3hMtEk1vF+IMOf//PjunsH97bUl23VSS1FLE3ssaos6RBCgTIxkaLiqG27loFQdOo
lyw7UHHzc2HnO3huojpobu5/tgBUflzC+sZQW9Xlb8BvVVN0lOSQDXUW0o4vdNNrS5uvHK+MGHvM
wErlcS114h5NFbHau1H5PiE0sGVLByzJDw6qto+3Cm6FpbpC0lHmG9v381B4iQxIndyaXRP35j75
WWvp3aSKAy3u8+kvA+xQKlNQ70zasyZ7sVRN5DAItJQu0lTgQHFYC1YlWMwXXAhstPNPhQv1VNLZ
jsdWGaV3owIUh8fgv+1O3s1EmLJH8umpSEkuwwTqQPyHGu4bvwUYfpkgc8BE93CGM/hu+lO2GPOv
2Fz7P+thkTfx2WygZIMGOmURgbIuq5OVoMU9dOU3F6X5omyVhthITxXPxIHKY04fUXx4vFMGNksF
RbBb4AMPxpPWZjUu6QdyfuaBcZcV9WlPLwXbnnh/1zpJiSPrsfXV1uYRqxIcF+WKnO2XhFXlNoyp
LzRVcSE89CNG8zTKBZ+NS87u78ZHBIXISBOSF6lFmgmCQZ3ZoM/djEZtG4UowccXMcORaFglw9j1
WpKK7TVnH9qzyJsvj1jPFQBMukqaJsFj1TLo2c/o9W08WMI/Gxx2b1hd6GlogY1To/WsfJv44Ob+
Uq08h/fQo0yZqFBr1s0qw2FSTUrgHKONORIFE4eoZsYkjcwGeZ5URZj3dLepCRO5rwlUBSdK8Vt7
uXmgUKtNAOeucPtDRSZZ9SNmad5M5zWLTjIvgxEnz8RCphm/J2BYPOu2/dZXgqVdoL10gqwAcRaK
JRg3EanzbtL80ShP5kI2+DSrEDPy/98N2yrlQW+wH101ApqeAJvx9V/noBsSIdQ/2jy2A1q+JLqT
x8vNH0otRouESuZGKrF2OArxJAGVA+hmjTeLL6uUk9DciXk/mkf1ot0WuKSgWX34fxT2ig9NoHa7
yNSrXwT1b1ogNvqnpo0x8nzgX770bB2rOjP4OmWjbzkpwPAY9+OjOJ08sABLt+zWf7S5e4IU13/7
4sMiKY34TwywKuJ8UvG1d6V5NmWBjqqgNOQKiHQbaphaXLYQDQ0oNRDvYWAObzqJWo08rhksdxiM
Gg7Nv/zRxQsP5mu94uefGHPzph7Y/Y52b3LJM1Em9YeiKhBy48uShhaYyYD01s5cGpnoGaVXxZv6
dRIYDsnPyK+73qnSp1IOqQ+mARKgecJTz7/1K8XmuIcV/FkJO2zd8HBD0HrfZUvNyZmYHcf4rRZs
ptHiYGuRUWJhwKnELyLx6Ar3VAKpshdH8iodHQB8d84KBCu24GSqynJPGwdO5AukCoWibz1kB+GT
oxPR9fFSw+m7ftxQq3dgQ/eOYc3+2DLwIF2RbhggEmrPkGRkbBSfjUtr8e44ze4Q3RO9ZuUdBkjp
C8dT6vP51po7vciLLrtKZVYNqWc/DXllXVK8rNwY0PalJ69/hTXkQcJ4sCfMcjQx0xzJl9uRT0fL
41+lMe2vNeOym8r2fglcTMeJJLfR+FSUn3oAXYzcokOUVnIgrAqgqeHRgzD4+fiybr67UXc6hlwh
SLGYGqLUb8RHtOiPBIpuktN11OVPAVqOGiGXVMfGkqrnck2XWYKHeuk1B8SM/256eEPzL4Zso/Lo
+UXKGky380Fta1mZhSblPpq6AAxmoEVy+yI8nKP4RloHjAX9kF9rxoqMh03ANInCoFWKy3AMbCfB
3BwwHLP0uOBhP7Tcaw7RpRolab2P9qqkllV8DgynqYIbOOV6cGO/A5VgzaIq48Q2h/6aXCUZ+70y
0v+5vQDRUuRyzc0q197GsxfH+Ept99taT0SXgkMcUrBdih+UbQO08Os9AX7hCN0WPUuzVNE/izUk
zhjGJLM9fVZDolvnkGvlTkQEfOVC2q4ph4CVEp2Y+sMQioiAcd9S5hAdT01wYBOQW6kcZnIJ2Hc2
zP/ftYJSiu697uv4ZeuL2m7kh0xtFa3hvPp3ISkCEmH43xag6uQN/6GDOjAPAQLLNWzeQNnRHDPY
TkQ6VI8xHcHtRgoTV8HU1zxpVmJJZk2OMIFaZiHTNvprj3lhDSa8p3atNU++liHjKVykQ4kXSp9G
C4uqfWTFMhvm1Tk7rKvFTpd3FeSMpvI5IjNxTiULNf+IsvAQKG2X72Fn76lRycQomXHCpn61HV7k
m9ui9+wrkvX5gsMsN1JhHkNqwQ2fMm62uOoCtKjQvmvW+ORbxolDP7CHb6tJyHRXAzJg2zpxLK+K
qILegidz+7YYWqAsNRj3q4RiMi3rzK+nEIs2CDnrklAmrcy3+k/OdpsmydUxYcDDwbj/Qqx1cfY7
O2y9zE/7t9oNSCVAzJC+Ravo3PsboOr9GgrfXpgQofXBqu+clJUJ/FJD+PfkYJzwSALBTkLTi3rf
6vObr/9KR3YVgBj4/CFs2bBAlnseMcZGpYMGkbs/zWmTNBQjuoT7rNSrky0zb5atwQXagUpulQga
iXm9I7jHDT6WfIc2O/wD/uXIRdB1hyZ93mTTolf88yDsaxi2bfcB2ysSB51t1zLPHre6jW3V+/Xv
Y5CcgzukJhSGD9yH7Z9O6U9O8cit0467pL9XW5ImuZSQV1iLVOjUbTGfkXMHMAeGsfiadEaezbns
CBPVMOKJ98TQYB93nEH8JWQZdILCp+HIT53Wtw0L/y+/CQQp2nuwBjCQpErDNbyN7gM0ojP2nnLI
Q/cyI6stWAb4ZrnQUTqNHY+z4K73OqYAgGQhqwVShlmTie2/d6s6v42SSsDNSuM/4nur2ycI0Su4
gAaJwaKCCDtxhJ7A2K3YwDwi5gAy5IHzkr1tmQ4emK/00YzT4WcbL6xjvOP9o+b1+e6MbWLQ72mJ
NZuay9DUpcK7Jxul/LXATMxepyUQOzc7mWloMut592vu5LbPfDeRPF338AlFi+1JqEPSb4cEQApT
HRkN7wyN5RJxLD0pCk2LMYT3TH6SSHm5YYFthUfikYx7QxteXAT8grLoGViLNZ39Kqk05uebaGYP
ptEEbtwzVTDdDndb77kYp4OS9Y5Gf43w4UJRJPsvCcibheWdqw33l633HYkK9x2LJOELVyPTRVcU
YrsyUeyp6MIgBjTFaruTNZCoW4KAr46V7gJ0+ES1Fb4Uu0Qx3PpnxMQ/F0XqZdVAsuhamK9Lp2Kg
flqQVbSHhx/1IO7YS1F3p6h27WvbR6WKSbNJFREv0JW2NtDdyA/zNZ3EHFxRzBb37axo36kiEHkX
qU05vfcWQHiHZgBwvMQlPOMQ78msBFMLW7AFHLyDiQrzNNkH1I6CQSC6DbyQXl/r06cS3UqsvTh8
+flLeLDfWHzq9wI6FmGuM2vhcVJz2rDwXTDzmXusRMnjwI3NK0rYWS52I8v46MjLNVWAOT/cAx71
0OtK4fzorczh+kiJwl2P9Fcrxp4SzJnnxfsHyOhFv39+daSowW3/L098qnnlQ+dl025lRxc9bSfj
ib/LYrVvgkLGAs8LJ3H3y43qv6z1PwbM+9gEeyNa4HzNPcmFLkjYAmf0M0mjid67CBatCg9RFc4/
SaK1V+aeiCVxgndScJ7jXWqfVu1fzUADwfrrQ/oGZTpECtJftBNARfCX08C7/eYhMz/H/MvkNDRY
8HPh9RWaJqV95Pul12aS6eKHJEFQp+AniUmZj54W8zZUTEMMqYT9K0MH6TfKmwHIIJpAqY77Ht85
aKTrplNnq4/OGnwFT9dWEHwDopdqlhS42003WZS4VELVBcjiopgKko0eaU+N0xRESo4x2djqK44U
XL4odRxQ2HNU1BtVDzUnDOFE9D1lzStjo7YISRJwcSXQ6gLcuWa5uRao9W4YIC1+rrCPJi7ZlzKl
cWHNOC0Fz5fEpYBfebbXCKZ8cjtD+mU4Ise5BwztvOA2EiE5NVtMdcK+I0Zl8EOq9yWzgebo294I
4mGJ2cEOyg70q4EHIghrESDj6MasKgquEh+TIjy3cC0fgw5W7XKOSrPA9d56hPlANHid2WtLeFGO
gMZNe30BpN1dlnnK9Uop3fk4ruJ2nZK4PBmH1PHxZSBrczkYbKEiZg6rKn0iDehxgEqBTsJLEGBs
vaEakVo4LOmb/JFE0+BmDjTIPHUJIUp6rv0q3O4cc+pCznlLaQVMUlr8eRw/gTigRsJNHTpSuJs/
E5eEUugxotGFDtrrE/N2rOaz5Se0JcYtUf9WwP+pPpVQleoMvHGQA+TD7Q4jTYiI8+bF+XDl2nFy
BLhSDzZEeLxrRdaijaoAu9uohknfiz7mfr6p1qUOetXLsnWdfbJ2h2NDpA+X2+3htyKGKqOC6++5
wenotRl+JRkMg8PHk1PRBRjCxk6iEUxfuF6TXg7BQ1asbiGv8oac4jgjxqexgeCZokEXFDakKVIU
o1yPFjXRwis07ypFGXYVm6sQKB/hA0OrDeDT7ZfrSX5ZC2cxgeWSfKZW5mJWgG2LzjJzuwRYV1eY
OuRDfKtH3xhaiQXX+w7XTi/ZrT4QLrxSESlnwIF61KiiXPy03OcQFVDqDY2Yof1F/RAE0SIGl4/J
BZY0KryXWjhOnWWhPn6aWI51wobfhvxrgAh+66ILmOvjVwKmW40Lq6ubeUClayuxEXoOyWle9wfc
PVpPl2B7XIjkMFusF+thQmI00nzZbuvmRfex5mlWe6eXXfCZe2jFP0VKdZMpdHpWmApiw6FLAr+J
HN3CjdUQx4bJpYBRChmT2jyCF9emc3WPKeYj2+vyLXZqv3i4ra7tOhGjV2QpSjDN+mDObOX1vzm5
VpFGB9ubPNHILlZfVlg4t9FohBGifzROPqNqfFjQ6kw9oKa1hjC+bwTTCIu+SlJLUnjJWMEak72r
zRqMrZIbifZlP7pelJaY01UDCjs953UhWD0a5HNSvgKftb7Ye+iSm1XuGqBNbWh9AUCrqc7H+6/c
CvwJ2mVdgPpdIzKfuUEA0Z+P96sTT1DEBIPQkEu+LMab93RYh+Zq2p+Vj9oV2HVZ/4olhOf1WtqT
NpnEanjWXNyuBtqIDGv2F4L6q/AkSqS6fTNM5n7NZQKphSY0Ux20uvJb1zqs5GNrSN9MI16CnIkM
V2M6lhbhOGyJNJ0BUWgs2jTVrKMaNdSz5p3uY3h7v9I21U+Z7XXm8xm59gk03dTjfEBTDuclyuaR
CNYYl5tO1xcvG6nZhh6E7Sne48uglVvNfMU6bBqQrYtwO63GKqSpR/b4FcDnaTCp7eBQ0ASfBESG
7qZ8N9lAC9NcYRpQ7NchOnYQs8b8qs0u+4fx5rAyTPYRYe5Wik014LkPjEj34fLqFLzuQZ06xLmA
0arzQUSRzAgmP9lZxySpzvyavf8VKcwn9Syo3DShOaOYxm3fcfDfgXADSjBaBb/owA8AyPVY8mwL
5Z+fWmM6A4rv6e0Buhqy6DFNMcGOfF7MwLT2Qvw43R+ALMDeOh+oS5ugM/vehLd9q6rG02RkyxuU
3gAwA87Tk8UThN0+dBiuFyRHCKpZSKZdTlyk8/7v3oTbw7kcBCjbNjvVTj5H8puLhSzBZYRrMWJx
89fofnkkDrs8fS6DBu9xByZDBDxXNiZGBmHwXmt3h/nu9AEwc7VU/k49oxTOTYdJzKZNa3/4Te0a
30PnZAiJRv8VBUnR6f6C5+nB9udpIwLIaLx69Lso4MdSFwraIffOgP8YJSNz32Mi0SElm7vEVAgI
9T8UPdNpie1SDUWgDwCBTYNBho0eHPe+KPCYVrc4Dt4LV/3l2nxhFYzxDXi6H0hcOxfuoh0w2Vqw
+qWFUkhduixRAcDtabaSZHbCDwQJZkBtJEq5cCmEvOVE2yGtaFm6UXHnqi3JleLj+nx1kWlZpFSS
gkEZipeTiasSd6cwzOYFxzNGMi+0H8AXpIKt0jOyN1RO1p2vl5C6PmtmQgQH5COBG2B6rKVtuoaR
YIwMcpuZLdcEtthx9an1LhnXNBXGyOaNUQumblgH4SdwwRXlstuklGuW0SGbyaIXLQxUE6KzStZY
7BuP0xl15ZArsVDTrfXHW4k8ubMyz56gH9vsPL4/H1fy6pyuOhkxZmuHkrDaqeiV3aaQfAViA7yn
8ATWlCkUHSO7Mbxyh8IMGnZXjn+PtgaAheikMaKlLb8oCheP3JGNGmresRja/q+zZ2tWuOOxXcYf
nhOONvOzTqgPRHvCRPj2zENEX55sIvQsZVzTrKqL7li9jPMR1P9NDtjeAejCtNh60dg+JoWJyVNv
zle4JsAmKloKGeol7zUfpWLQxcA6dXaAy3kt0nT29aUyjt2cLS3BylVGlsMURhZvp3nDD/9rSmOw
H/OdQHT+nRt+iBuzoEhpsAuDbRNTJz9S5nwNRTKYZApXWWByT+7A4sUTzB7HAo+TEP+ET/ZKnqY1
h5qDCfSpp7MiBmQfuBCCVevs6+wrv/77XqdUS3MGQg5TDJhyl3mh5v28EvH4GfPvvjFEnWPHpGKA
XV3DjKu0JhY3541Ac6p4L2mUnYOC9NFguZdSXz7sNZWBrwz7OKvT77YO2v8x60OnbwpJLSNvgW8e
GhhQ+VjyibPrgSkidm1UNnxuYUVTBxTN3iwRNmRGVtQqnp8exj8rPrno1f4IKds4ruZkxwat03nQ
4EBg8zO/DM30AM36av9wl9i0VcedCfLG0wDfzJ6Tvjqo4X/AUV2C10cCKDXP4THh+gByWy5OPcVd
WveKjrcL5MXaU/f5fUalINK+qsHo2KC0cA7oweIGLetugtjWV5atUFuy1ZziR4T3geIt20RlMqG3
jdyJtbXJv4cATDlpyMHFGl8m8W2e36/GcL6LE9dg5YY2nOatpexHkYATNwmYebtMrc4GBzzxYFgc
I46aG1xHkpvSRna0BHWapY7TEr/e3mBlcdjW/dTS8I0NAwHrHMMe4buIzKXOjTKz825AOP3FnrNJ
UHgqGDG330Chmt1lCgII+mcS2fYsSMYaBVWVlT2VsbvyZIPWpg8DzKFEh7Olb8Vk846aMOqoAkSZ
IPpIbjLDNyfFjFmjekrVv+8ZfAdE1ZkcTKVa5vAcJ/KZVWogdKSl2fiMs4IB5vatrWx/RAClACT+
JQWN+2DYxThg1iRJCxrxN0A2Dv8wOJK4UH6gd8ICCC/SssJQdQP9DlkvW+ERwTfJjKAzGaJud9E2
jHoWVAUm+Z8DdGjNmrccxR5sziqw4KtnKgFdM6QJ0RA2ocYQRUJgg6ZGIa0UKNDvcOLS7cM+4EU+
wIWjRZwQxyQ8vGodGrT4EXIgLDMpBx8gCJLtkHGti6kKT1vRt4kHsr6jAd0tOklfNCxzm01+2C20
09a9FzDEQ7FvRbsLc2vJyKyE/xhzW3+cpQ6GHu1fDOKxDNqn0EpYbbAhV0dt4SKi/PF2kf6540ND
T4qtXUXnvSc5lxKQ7TKH2/qmbvLkxU1yeVZTW8Hewr1dgmFQcxyGrJbwvyYd/wb+GgYFxCSHBgEB
xi+T9utDPaUj5CTRpuGjB3ui3obcUdDjK660Y/kLqGqfZEvtND8pZhjXjNFNacF2/yzO/JLPui9r
eFDglBQknpfFymYgrHOLwNw3MYNGPjOIRh5Kpk7XSDUrtmjIYKHL2Q2HMCvTMyZJqHWC0AGzhkXA
zlh20AX6tF4lbTo1eUuB4r79J05YLFdUjmBNHHzd0pB3UjweNOssMmgxWaeEx8qdRdyIVQtdpbsx
FKTmAQ4+TvXHunddWZGSYZv3NTIvpy3JRBNkwaaRRJQCr4TicHxOfQrTQLDpbwEfgan8UEAkoIvM
gf5AIjhe9veieL8d4Qe4athRR5L8Wst80kd7nxAckENQIWpfX02plFeiYQMgvHMA9ocK3/Lt19Zo
RFgXBNx8EaXazasLec413qflNXVz82Ksge2W92W9ye4xulxZ/xajZc190icBMLR+V00SOD/95j3E
n2lr2pvKHSsEgRNmuRPzbVSEt6tgRG0bGhFI8sHx0mF8fgb4fbuZ0lh5taZ/KDqS/E1aA/N16w4i
AODtix6qn2DyIfO2YiImmhvWZ+QcAY5MOrghN/4MglwCiD9UGHwE07KRAjO8iNNXiwnQvvXlZpZB
Q/LmJht+zPthK4HR+igh0rJ2tYPD6kVqaAEpyMar5lJdoLig/yrREJinE2IcfCUpYLHR7svRD+MH
OS0KPnoufUsWR7GpKwlOA62iTUcUvHFN2LjLuE5g1m3EOI4x4hapavTtMpQMJtIBF8N0CFR1wiwX
2lplOf3p49QV7+9Nq2kPS3ARfvtrh604wZF9fUaMczel2uTQ7j4hFfC0RmeMK2s0F2jUzOOkWHG3
Tq/7CR3IsDUSkCWU0WnP2peW1W++PtrNj6dUDjqVRDFS8lDFiVTxrSK9om1di4BlC/wJ9GCIFySL
rVc4nJg+J00LMTRX8bQZ/2Ti/QM7iD7GRtK6BgRrhWamqK5P1SsX3qNYAyB4pDNpXYQZv2ljI3Jx
TmL0xcw70iDDdKpxoN7voJqjYQDgjl/ZJXTePL/HjLjFLmhAyUXW7UV3UBQsbXTOWmB+aNwt3fnb
LgVY6soRChYqMrqT/I7YYboPfridjoZpOR61KUJffVRvkW+WWpedXgpwL2CgoRu4RgCxU2VdYqAE
mWinYKhrLLixpF9jU84x4WWdtpZphV2fC6GYvZAZtldgC+9gQhAQ4kxBDitjlhLPxluhvpRiM2d2
s1MtIx2MXFqQ/+EVngKCs1/dQaWNOnugwC1vNPA9ExPVil+wWWuXsplC0Bt0Bdfr42MGMS67+vXH
2U9RX3zUm/dcVFUhdCiAWf/m98Wt+pEsIXkbR5gQC1FinBAHIjzswTP+69bKbu78ZV34CJ+Xqd6m
NbPGWolTh7wdBIpkYTWimju/KUvSA5WJgWzJcKUn1lfTCtZ75hZxL6wnRLz/A2YIPdONHwHAGhkw
74/9hF7/5WT9vdP853tin/KQnBlJb04Ph/lk3yrZ/MNodrBnVvIQrCYLSdRNHni+PgNjtuQa9wIH
tTebPFd7b+9pW+Y2B81vKzVLyJIjjARcgSgW4GwGxfnPOxA9BCh3FuuPEwenGlkJly9cWxRP2jKy
M33A0eUmVh3NggA6LE+pVM6yzZkWVTF0CwrTc9kKkedRryhNErJnFdYnpuFzIH4IwuV89TpCL2Sr
9qyjgUL1xWAI5kz4834dJsosqwRg33OVTJIhAJkR+1dQEvi0YqCBqx4AWHQBRYP8kj3sisMzXSgj
m/fnQfGi8WPDqouDvEhFqdQ0i56uPgulo9qP05wGcJEud1ICbUOhAjnEi6urZwyN2sOK9RZKRCoh
oVHYQAXGCOY4YRRNMZ3EzIgTmvj1KDtgaZptV1RKOVE8EkbZRgtNOV/3YWtnlIhA8EAViPPBXrcC
bO6GZZLBrS7Tx7XzaHz7zqn84dnavhP/E4tT5mmJ0cQlojOFA6QRNyHt2qG/cJcEwEwlYjeEOSEB
AqJoaEqQuqQ9O94ElMtzGsE8FqV1tnUnatEvEv8gPjGk95ymXi17PQDJp+OLd8NguJNKDsaGi6IA
iyudUuf54UE5tnTgefZT0qhyzPK39LivtuZw/Nea6wS+Sfpi1RA0qG7H+xZyQ9bpvqu+roFZFmgU
xOpUshHgX6seE7ep92Q68uyxK1vHw8qGpjFEjHW8FTKRp1LwibdTsYntdbitxoN16AWWwlmhgyaO
hUn+DZbi3MsA300N6Ue1dmZLo2im2I6bCBjrjBjMbn2UE7XNd+LGA0HtMoFuSgDcU5tAuyTVE8BT
efzA9WsFNMJEkCuY01hSc8aN/Tk3rgdT9Y8G1/Qe7U/eHMt2wUlK7UDd3ibL2mYgGyikawWKGPyT
2UTHi3Is3hfBB6oSm7b9/Ix0ycYIxk1iziWXGEDI/aJcE342bwTo9qD8A5wtaBx90DHgLVcj79le
TTUQyeN6sy42kBs5NWnfAAmlhdPcPoZ+O5B2JpV8lVAkSbmarCCFG/Dgf4nhrXApPNATI5xmr7ls
kD8YRPSWfG5ocWjIwBeth0qmg+2MxLsJHL4BGJTzrfh/XxSCJ58tTSMZ+UfncPvfx7x4VI0iwiU3
c1yh7FpjPD3IqGVd5xAi/9sETUqhj830pJHE7FO0vy4Lytd1EY0ARw3JKSsbcl9H+LR+DTrnreIj
UhEl0hPzFoubSlp4X/tdyqNoCbDkDd6fDGLEyaaeGDhgr2v1d7LuM0gG9+qORHfC0VbCwMG1YKyC
xXAlDldivu/5VBGKG31PQvlNcDppaRFIlDxpTYsw3EvAF5acq2PK+GrfC2u/y0EVFCE6LgeBariJ
hwVoX+Uabge2UKiWSDvrtl66LeToGg8hseEn0oCYMVxu8uJiFGmSpgQYSN512kl77SXJyblje4rQ
bVtdFIMWVdHpiP4ke4I2FQGzkdv7MjsAU/U6td1gjecIT/n53dolaH5gGPH1UZE8NkTKPPkUB2eP
yiyZrG7NtX/wrvvI3LrWqVhf+9f+Y27GeEpmn6mKkgScfKNP0GFVTuXLQUkWOMfunbcRKdG5TSqb
So8CQJrLB44lP00qb1kxNixWOxvPVPaBGVyWK3JuhGcmamPFV0HOTTnLeJGMYnsPKzTMgMyHrFdX
mjIKLf+VWzwci3xSoerszn9HBHxpYrBsNQtySN5lK0n9fgiddX4TMWtYs4rssTg/Do6PTbbtzMTr
52kOHx82EQWD5Hwe5N7kNDld7xJkARsHWRSegAGd1U4Gqp9SNkNqvxKmoJL05HwNJdw69dQlG8Pz
FZizJehX3FpBSQz6qkVRJlbCW3nhLcaau6nEyl0EqAtTRrq8B9fNobVSw7L5aZdisBgGkoplChNh
n2uVk/r1PmfQpfTlZ++dOHsKB3S5hem364pNCV5YnZSZOgPCkE3rh8rcsNujlwUeoCbkKmxhHg/5
N2Cg9io4NBk+7wCfhyQ8BYZR0tlVPgXd0cFafKrwDdSkRlNhYPlRjeCkJ6bAtgyuhfkMnsgo/NPE
hB3M6Pw96BRpUHqKpP3m8r5bJci+bTrkmAZPqfmhPHqvJy5kVkzXk5HpsAC4rJEIJSXVfEFXT/yi
phYSNMSQqGdOG+RBmjRAQQDjeLXtOLmsOCgKoJROeg+UvmbHbVERUzXZhQy+ealFZFTXNrRq4CZj
J2kqY0ivEjGuarJ5noxFqSrKr8gHhYzTmXFY2iE+szOrJYKU08fW7U77Pz3KXAtQ9WYTRQfvWVGt
7OCFYcIjBFOa2opcnvKdBRyFp3jDTKud50Zod17EE656uyOVDP6RY+/4rXv34Y7UXuu5DBWWAcI1
AjRIROjKgJQI88uy+HsnMnxWukzd+QShXFs4NcqEPN7j/SrN+An77mdJFfqoK9LDyLOR33m9P7cL
BlkvSZbmVQypbAUBkPMA+PMOzsE4526yzhzU509mPiuY331BZE3Kja03SERKYgSTv8GKK45mg12O
hjMbmwZRQSyL0WF8FT81vb1MFfApK+gKb049xmnYCaCk6wxPLv56qwwQbl1nTrfjk+mmdDtQ/HwF
2iy+zBL4xmI6/tGRFlF8FvmvcVU1TFELxmDpVIGQZNbLR4sSuoyf5v4VmptYRQjrk/90IM1vRftU
Z8I8yjECJzYFKya3a4y66Tkl+oUVIlXkcxhr2sIX8aiMDK+zkInZL1EbbfGx/lBDFeNYjQW8lOYa
HYmDlbkxrKmHNMmbduU9hRaLnr7rfJxLJr4N1DyBAcMMH0E1p1ipsmWSqH65gEbGye1beYDTPEAE
PBT/xNAzXO2QHUTbMaOtRGUbj3Tv91jFeWtmo/LXgUDVE6muaEmp5qiYkj+vVU1EdUhR/D3oAzKD
p+AU/NmucnxF2DDuNOclEL4bWvk6rFc445GzF9v4W6C1u6cYytHa0OA3EPFudSn0o9lENGtLE2A1
uqNN9XO61yucTkDbia8FHfe8gKOngOdT27LQ8/ddZ397laDt+Yp8IZ2V4b3l62Sov1gY4OW5LcIy
mLOqnfh9k5l/WafpROvaGk6kjbLCP5f55WHog36yCweyjITEENL5e7KTC6sw5BNrLdWoZWGtPWRT
S7+64Xixv7wad+Q6R/52zUUiE60FbBpubd3kM63WeP4fGsf5vhhKvPX/vP+awnFmUqvPVcWSZObB
Y3LCbl/HHyXgcrGEfm0nkRZIzSe8EDlahTzlEdFUNMyrFYj4B9b0WiPt+3u7+Tsrz7cB8IECBL0f
ZUfldT3IQck07ASkxBlcNE/1z8yKkGKJ5MyVp9sPzCAJbGWFJg23+bwG+RhJWFt2AEGK+nZpL9bw
OBZloHsllgCXsXhu6MWgDHad4cYP2yaYii1SyENL9Npjk6RzLpS/ksx5mIOH1r1v42pNPzkIKZ6e
mNcVPxgSRJm1esWAY0gHu5imZAKvK81k4aQGt3k62K+AQ4YHqO/3KYUW+h8C0CeUSD+RkqzCDs6S
/GiWgcYN1E4YLcS9LunzsaZBpVv/mOhcGBUpcrXYI6UlK+4gHwEVhatTQNoxoOvI7cDJpKE+UdO2
zbBAYd/y3nUq1Wd8TSm7HX5hhSVXk+4X43WqpJRLBiGWCluwrCNsNwGM2Q4X9HXRno2ZnYM8eL7E
X4SP8AJbiKWO8BpzK8yg81agoJk8DZbguJO6drMaElustoRtl3on6QIX0NTVosp99mbTNPowXggr
/zMdj1Sjc0yDnK7TmvtKo131/s076Gn5ytpGuKn/dQmfWNfAvwZ8J29yq7DTeirKSo7jSXjsrNSs
tNN9PHCPIgv+fomegsU10sTHAPVXOVoaS8R3z2KxTWdf6eDq2yrKGEfpz6F365BzshiIunACPLRl
PYXG9WunNct2FItvWNSFD6Rg9dyej2bEVlyTPt+ZaUVHtAQQD27EZdUtM43DE4IoSUDVKS2Un3KA
1Y41bz64iRK0knAfB4IceNc9AVZzD4pt97r8h6UUp0bK1wsPH6DZAMGlrVqtk06bZsdDFHbDHKtX
k14mvU9/BIRvzMmSQZMyZHfwkvRVGYx2BR9IChgnymyUd+5MR8+JYbCkJmh6C6hKT6mN3wN/oZSD
SyAR7cvRvQr3/GVcIcIEBUVkcBUf3Z8b+IuhwO0Zzby/0sxy3nSn5wh2TPglyp94NcwJPlkgL4oO
YlF/Vh24a/6ZHGVOgdhQOVZAKTvxT+IyYx+hKFZjrsNE/Aj9McYTQyK+jGcDUMc88tiJFK1fyTN/
0xyJQ5MtAuIfPgBJHLZGoF95FUKorBTWJZllosGCEAS97YaIf/XI2DlwCZwTZKpOxByIiSDzAgAq
uiXwOp3VGYxh/vtJDOtCc5x8WtYjUp37uEjtoZqfwKPZBH6diSv37gU+qPsJpf7POqhesQUnaVi1
FTwWcUad0E/cT+5gPOLOSEKouSBH39tYMR4EEqyMZ4SDpRP7I8Mg7V+kLJkSzticsZ807sRfUSOs
B4E1xUJW2HXvaqmCR78gW8spXDjRp6X4bGGeck9A9vF+tgU68e/y0EIFV4BKZfnXbLJknGHvfuJM
p3tWVQ5ieIUebXBVmEopniIHUCjR5bW7ZXOTK9wXiR9EhCNMqBPL8vMF9msuamw8VuykbFrOeGV0
lGvx8NNF5IPKkMpVfCqUI+o1kWGJUGtJD/qalN+nmq1++6+Sxea4V2XAwBaDXSXe9XYYgDd7WZl5
QSYPYEPWhO45Qj4frcJagwOi5JJwL3DQ+TpVPYMwFf8Dr/+cG99KCSGCMpZGLOo6Tv7y6ZezWh4j
Nb+lwoPMm9gJ9ZH5usVIuWGdAO2lGgZkgBzECk/F+PDynhWLEfMzZN4D7iHIEPCRS7nXhrLTtkSO
sFUoe1zlsTf5zZQN3jF2wWZCIKZOxx4RPwv4dk/S6RK5OlYSz7cnEmUjMTA0JzucZuC4tjtZL35J
RF1AwZ0AaFH1FmeUZBDZdQx4Fp5qwCXLB2X7uOesMvU30kk8aYjcT3EoXAesNn3TCeyS8/oFmNts
cjCvLUPMSzm/qHj1R0oaCbLcudC4FS0BjJ6rPUAXa1MqB38l9J+Kio4B9jTi61qrenvy8d1b1TBB
0AGvX8zWpJ6GHRaMXbS51Gj0hinJPFhEcQLSc+jFsQC77Li7IUs+5jv3Q9UURt+qnGHNS7BV+C26
2nJZjgQCUpG3xZd4BEHfHtXXYCFO3IG7PBuuakemTd3VLwmEmHZkaKakvYDvemUpN3O5juEp4d31
WxKWmpgoPazDO4Iq3cPcnBElIEaxjDXhc8uNXP50ue6/sYEiu+6VIMnMhSS2IvUFurtytAmBW1nO
/4V1g/n/RVdgaeTnGZkjpWxmnn5cMiiiN9Hw4EqQqjWKJ2QAxmBFHrJHpC80OMGev7ZmRNInM8nG
j8a9RqMhh7PQaoNR4MlsUggqZKpk+iFy3zm0rBqbryE3gDmvyZ4++wGYtk5cKegzP6bRipyeaKqx
ktDZMIi2ROozS0WzztmMKXAliJ/2rIGjxyf5zS6d2T6I2afTo5YB8va0qSwWxo7X5YgS5YWtXrde
hzETjAGG5hx+od499TzsrW+EZFjCIQ4BpJP7m2ZifHV6LkvyPaH0fi9C55XSJEtlGyOloMfbaIJL
Kg11xIWf3y2JQkVf1MTq4Okpr9LZ2bgUZ4k28duOdA5D5rRvJPMm49bXXBc9x70lhQsJDFwgXTRY
7e8V/gxRVTP2MxF/qdan25Zl3mbj/I5iM8fSLzLQAit+rm+52mkE956fpU59h+/nLNUYyfF3ygMB
pwTwCH2iSgPcXOFglTc1CmhA+aeeX755dWOPjL1OMzBghOWdO3j1L60ws70RzMov5QZ+9zMKPvSN
wFjbVeUhW/FgKOBLnw0OXPfjqZ8Nt7/38/389AUbW8aUl5Ndp+oW4B/KpTQl2Jf6Eh3ws7SN0nT7
l764vFe8u2LJZKPvxyOrJfzAayhw6KLz64Yt1+AfSQDC19VfThJBDpxfeFUAKddAudZ6Qb3PNUvN
76kAO79M2s3T4ljRnRY52FkoBu9InpKIKTb+XUYMUBo39EMNqAs3pBdEMYr29zfaXFyU7oEwghj9
YRA9nejk1a3QscgIvUPpLvRYzwFpU+YLD/vdjdr+rSVA4fCpxlh9zTgA/ifEOyOVt4EArR3uaXSe
vVTvLlHnwvAZrBxz96wcwZgys1SoFtRCP5McAtq1xnS6sA9oK5iQto8JggGEkGARxfmBStjCUkte
Rxf4pmG5lYNO/0uNxlvs8MQgcpmDQhisy+DbeRhQnxmy043JJtcFZVn7hyq6kEAgvbLtTTpNVXM+
JZPKzCiSdNrCbwwJfBFv51BBP3MLM4fSZYhuBk00jiM7EgjpJV90SsG3Ojgoh51I15hCmAGfpqxJ
yMv44LCkKF8vIjWSUmpbu96Jub3BNs4FsXxSg2feAIs+LF1KxKumN9SpIbF9jUIAqVtluDvojKPc
XG5Fm1QACvfZD7gCSRuI6bDlsenvtL/4O2xp7Q01scxI3fFNxY2WwHwGzRSGkXLPiP1hS2BPFyel
5znj5u98xBHnhoQGHbZZ+oTu6e+Pr6Kxi/CwqMwJP+CRmqStGnxCo5HBLdZC/ts2A0ZfvveNQWJ5
eaGaT6DRyL2NMFtXcnB/yn82+DIRY/17VB4M5gr5uVlnH0qxvTWznaOaWmiwT31DkB9E2Mq1FZaM
f4sVYHAuCqZdcZrXH/ee4bSsMgF1gfGCFzRAESofE52S24D9GD7NwJz+rGT5800wi1pG/1Ao8PR3
FdOU0dxj1Jo5b+ZmTya8Ct6RRD+ukyaNeuhl/A6SaPRnZ9hpnwbgO6ZG1aT93Yfl9IKvAHE9s9jA
1btibmJ0yiqHdRsJcNX5wuZeVdEcBXE78wZNhs+/GtvrOj1TZfm0fQ2peMfRYp9GOuRwdlX+zQY3
OwGJhbTsgMLgz37intcNIZVcSgzJotJcR0OWwmL6KEVMtTpjxtb4e2XNMytkCY4LFRrZRW98IoVj
Gq4vtlcbuierSpXdtW17coSG+TrROCsXy/jqAaH++bfnDk1adheLITyFlU8qCXO797m09IxHLTof
eWYC0dfSiXicwoCbhpTrUbhMqLOP0pYkcVDbgphLnlGAWfr/VROngk3KEf4mm4/sqvorBHYM74vX
7I0bQdIZqPWHvirEIyOkj9U9mtK/T0C2B70UOmyrTkyc9cpXFtt/u6/yYCBSGln/EmMl4XY0bVXj
sRAeKByOVYudUIRT6okeCbHU+C3wBjimf634n2cqAQM2XRHL8FulkYtIeVnWwBpgUFF32E0k2Ize
X38iRViYyUtaujWd5UkH7xUL5bBpb2FDHQKnVHx51ZLE/yUkKCVqlXv+yypIIqK4p/bit8nuqg6r
RU5xpHLSufaYFbkl+jjcIEnBCSu5MVf/srxRPucfCp2cMCuaLx9qQAczn8lw81Ks/C6HNpes2CMo
VQ7nz1KEeqRnViIeNwxbvSY+WwtPTC1DgNpKrp86O+bpKorazNP6CxAyAEVya7DBm2zsmaHHm2Rr
4e+EAu7sUTZvNrYP+nXNFZFrDeE9QHYnqcfrF4DINSNYULIB6MGP4iDrKFE1/REM7QVSunB8GqEz
6VqNgIUbqZZArTVuVTnjKcoFf9ArCG9js8lPkvUQhErP3ZahvOTxEAqCd+8luVjBX4N8LY6Iqj4b
3poP46QyJWTP5UdHOfbDM1rdP4TBBBFbV0U1EPwn61E5x0UWUcpqGUEnjLzGqLYbItUEzeK32MNp
fHhGvyWb0hoL6G1BleJGRzKJKQgwyFSAg8WvNQBjuLfkhHMpWw0GKXdcz1z4eVYaMh3JTcvkvJvI
xspnFylXTlrjrYd8CQIf1YhQ9vxp/AfDS0sVBij1IkPb3YmYcwLu6I4DnuHcarjF2PgRpb8aNEdv
q+6oHSTj2YZkYTGZq5nCbONNcq1FUB6PbfFr3pv1tXI5L54MhfblqjvRL7JqaT7xiTTdrl4Et07H
Fo7JBVnnKd3TyvSDgjkrzzUp3dulQdbYQT0udHRuk/90iTOip8M3jfiEMWodSDuBcLWZ3f0OUeGE
/u6lprS03dyi87O1xfFtdvBjZcfwLC/m3Sq0kbv7PHWfv+PnfGmtCk5da7y8lTy0yyBEakGOWhp2
5lVwh17ivJ7fphxQ3YjSsktP2A/KcVZPN1t2CL7J2H1g0dJhu8nKoeI7/s7xMzIY8OBZLTjGZ56P
vl0QwXe/mTALVdtf3ZFTbJnERL5F6j326wZc74dkPagz7falEsOxK1gkBXCyiXl5saTcZspAyGJp
Ci5+tNrpwzIMQAnc7f3ucXy1AvokV13BqRfcl1ATtTz2zyXX9oJUkLeTYWIz0CrVDSFHeQjcf1f4
youL/URG0gtEf5ZIBvhvHoQpkBn3/W8S5kJJaanu4T+5IPKcYWKicRW/P5oKUwoisVzMWxWPlJm/
h1RFH6hrZaWT5UW6KUT1oA764vgZkLC4GU+mhF4p6RMRXxhdvjJkTrclmTeSHLbvvWQmXa4dnW0e
+oW9yTSkl5uyyhwBhx+k5ou85EwHu0S8EczpPysZYhD2rn+YzJMYrpRtqkVCf8ORpwjArj7RvDEb
s0qs2FIkD9YUffKzBKsFqYFk+J4Qa5HV6ffRIEeDdqDHH5gtKz6arCwrWRvvqPn5dnC7O0bI7hP1
wYJdsnqTv9InjLnD+RjCLYVUg65KygSICVB9CPjygjeLPsr2tZaE+KYY0tECRpo8G8KfGtmsKbD9
dtXG7htyVOW80gWAAOM7eYMVNU2UiwGHK59VBFnerZljune8+Qk8CVDfUpBE7Scd4zRcAXNAfYtz
om+7/9dgpMTYD2ApdvpXPyOk8LxeoyEadDWOIpP7BRDdATeDvUzGRliK4WgEYB/dJVrG5nBZl1yg
E4JT5KNjsqHoXTdEiGBmxKJihH4MFcGYE9gRCLqNPvHTtrsTuAvE23hj2I+ZL0CZobYCEx/MoaX0
mx+42059UERiaA2ZmszLjH8bXeOssloYVu7/Tblz64H2sL8shFl2FYp8eEtURP4IiQc3gCLrkDBa
sSGuBLCUZTorY9imeHk1yJvF8qSGRAXxp6UBZDW/JBPYU+cvrHFE99ctnl5cu+Y9ZXsnopehOrF/
gUlX3MvpxXfja4/+YisXOlmZtAH9KWXSFli+APrHN51OEyppCg3mUgQWfDettDRllY0v2yOYGgi7
i62sc2lEE5tTdEdLJtUvXoqaGaeCxE4H6K4EwBAwIEcFFYHHONEDeBjr5EdDZi02m1zx+7iFpgZs
5t6ZE/u9hH4hDneY7EP/yMREWdwxAwn62PUqSQBMHXxGRd6naq1RzP/kZ68LGxfBdvDLXoaEE2v8
Tn3/SIYlaC5nEm6bXn7FJKrJzhX4TCmfDXGA2w6+tbqvsnPM5JTUIWxA+lmREiaeGd6tiWb7c5hZ
lv5SVkrVffGMKzSYQjmv8dAV57aIW4fHH/IjzsKIBDGtAKbr0rfyG7VA81+c+jWp/uYqAmnqUpL5
Qxy/+TGo4EkTsNj8L1iMa2r/SuAMQrB97iAaEahV1ZQ0RZ+uo3uzZ+gwwOqHLlD4lK1p4MfqGj3C
yXnXO4Ks7ISbkSAjxVFgM76oAaTA0zGkcFYbM/WKedl90dm1YY2+ANY3OhX8thQeuO8EDEKuFUQO
LLaoqAo7kOrd/ub4eWeUwwXWYvV2JYrgnhgFCVdrnxesfTEOB1ubcJPH7+HrWXODZyI0qU/oZHmF
Wthqjm6Jn2ZmMxs/ObvjGGcskhknWb2wKQELRZmpExcEc0V8faNK68lQkN8sOI6agUpORlz6Airc
Y7h1e0DMP0dJHeiauWNyoW70smY+y47SdY1pyXspwEHsRxmpOOKqfjYNVsy94eauZ8j4JyWyY6Sh
sAqAPRiiTvfVMQbqIPDqtfqh5sMS94wUzAuTw4sTRYYFe6AXCXp8VOOX8YdAXwmw9iH3SHIsGpYq
546XEKoft9sdXXNT3hekOVy5vALGSuS/T7XuosiO6z+lg739PZnyFSBaDTeEQLfVn/6ERu0bRHkB
zerrkbQFIJttWKXPpNdBn7ZJ5W2F1hkaTqPH1Yoj0EjLIda+COFzHiRvzl52/PH9v0DBl7wbHNro
oLdVIRJpuGf+hXK3gHG5ZEghFjwPQxRRMQ1Ro1QRwQ8Du7PkxsEk1TxnrCSNZ9AuDtMlff0eNxmN
5rhW3vBFbDo5F8q/BVKVX3WLX+QTykKQP3pt7iLm837j80d6I7GaHnS1j+dE7XtdMs/dD51wmSKz
Tcj5HLrNOnCiZY+xLjvvoAdOxgGQprvX48WPBe4DbknGiaZYJ291y6TTiLeIl9LDjlMIXt0psw28
/kw9W/ptO9qMfrvJZOjTGRGdYzQ2XdnWMalFyisBKpHKeuDV4yoZQJEZbzDuyD9/5a0kusn0S0RA
SuHekZGWhPt4yXerv/eTglVFKxG9hPik3/riEE5yREOtRFiu7rfTKdmSp3Dq6kWW1U3eW8VRC1dn
fV+LDoICSQo+F32PazkLYExlkvaC8uJ+/AFXBdZXtAQfB9HF9q3rve/1X0PgWwU7XIap4e7e31FP
+5sfjyQkb0KhctgSbwM7wXg5uv/YmZ89IfjT3gX5hVHtZ+cKBGUBG7f6XUBGWAjV+rGejiGKgYv6
Uh3m1xVte5YZ7mUmxpCqYIdw+yFvO5mslt0qkQtHjcTnFmyJvbPriVfROb6A8YOscuiKzPz+/2NV
St1c9QwzPgXozrGSffMsLm2z3uh9B7v73txfhPdxopsf6HmfI5NWlQ045nxSP3dZ9pud6B/JKrqh
ptFXJX6BABv9saW9hmE8mEdmD3zUYTOoVaR8wGx5rEct3ABLD36OapYt9nQjo6t1UAYWED1xSruR
f1ACo3pdA3LtwRwKp+zfVs3ky/vDhFm/TNk4jqwzWEnf44llY1ZGcrXa25LxWkcqdVanqosQVQeJ
C2oy+/KJ9kIxsXkz33vVCKp/Yriu8Rb50ifwTtgj0l3RFKfICyXFg6oE6lcoDKdIjMAsdrLzQYeB
CPU62ylkGAkn4HEVMrztuChZi7Gxay2M8Im1AYZFKjA6pifTfR0YORYFc2nqtxwGKsmyM40yldUU
qzkv32WEauwmAqf3+MFYPKoO+iR3skvbykiXrJCTF/ieVHQANir8NTxsYI5kCyvmBByFnsAwG0Lm
ukAqmmiMu7ZkOr7qW5DvanJLc4ZeqYEJ65bEUYkWmfOFHdq16DOjG5CnvwSuBjqyThWIZjBWvhRU
zID9Z0PqfrefuF3kT7x7epzw4vc9AFutnOofcx1+QTYOPle7vT4rHcRUpmFR4EOnevixGnWfV4HQ
u5doK8x+F7xpv3Rkxnnsdoy6sKdai/JePI0L0ijaR1RusWuA6DYOYY4ndV1iEGn+rhdG9qaFmJfD
cFnfSAjXjxDnuQIbH5AZ7sbTV5H8fEoSIZpsYWb0VXXRKjpNdFMS9b3jkEnh1viO4hfhvT5R9dDk
kLftelW6+DxYVWUQS9xNCcs6Z2dJvreeMYuN831x8w0hF3C2J0Cxoc27yn5QloGBeSO2z6d2kbO6
RRuptat4CRWvAtq4AJbuCahDz3NkXfgz1bvREz/GkvN6qdLG3xU4BnfosSQB2xRw9GSuqFNjkXk3
jLt9ns1St9KfuW0ZdDJS4XCXp93SOS6wjlNqKgIJR9TjOm9iFqP9OFyCnFhU3Ep1Bv2wEZjMDFk6
A2b85x2I5A2imN8Ah+nO4pdYNB/CccUmAP2YBCsoDMAulCeT2+dnfsekxhboMF6yG8zq7+VQv2mo
wZuyhvgQZZ03PHkZqHEP/8BKpfbCeydABhzCPSHaW+dr+6beAJ+tkUw3zPc5oGmzvVK0C6gfU+vA
CsKtXV0y4/I1OGKFMc6uKKy38ETQt4fMUcUQOUMBxNlrOgiLCkTh5V5InReEeQKW3XufOep4HK42
REdzaiTZYJ1FjSwz8EGzzu28vh2vlhTCJOZDN8k8grK1qQHokcxW8WNSdlay9fo2YpJ83uJfwlj+
XH/++R0/MfiPZ4zyX/aDWZGifOEmtF7KT2eRNt05KIJ24uMe3PHceLSUjUVOHKMtVlrYHqGZjwsX
22PyPPFWem69jypp2UG+arTABcr7FKCcrRQn4P4CmfOM7JUzmV6odzIH9x3wWMJjNLfiLd5xumuQ
w+IDfVVgyr4SUPxPXDzQAEm+ShCTac8671Y8lPq8JAmFlju7xUXnE2PpHLQdoiCoLXYfEIdl9fRH
Z03UUaIeU9xOJMSUVjbUydEW0ptLoi3PqYjJy3KbvFF9F1PMhdni2h8aDhI33C3qnnUhOCXiq1+m
jKIl+gEx6X7LoGIOOKrhn7sroiX5v7Ph1M/4nH3AMzp9SkhfdOrIpH7BigoUaE6JPyh6HH4SItwQ
guAga9cTPzSt0qZTAYNtdTzw1LsSVu4OTQDlcxTN26Y+EwOp1Z2Chyyrd3OCKTcufRxJnlkxMDgQ
9dlgatA1QPcQUb88j7EHJ0Q8JDus5SSyuwy4bj2NLNX0zs1NBBYAmY6kSf4qDh5GhZcTgmWqbB3r
tPNGdQieoNOaU4uZKvB9ye9hQyTJQnOAqD/sFrcYwNxjYEiVyM6mK63TVOjvRt2PQ5fM174dhNqZ
aSfWdi6Cb5gFGd6Lnsw5pXl+8wv39fvOn4P4IK6WvW8VL2fyPatj4/0D0F+9wXH4/i4528zdoUAF
hT0o0sxK5zBbMx7oGa4CmjIZpoPZ1fadvsbmyI2c49MWivMYWjhBjFYatgc0x1hVc11iCYuooLgV
qhzI/Ad/6s2S8nqI3ZBNix6DR9gLv/oYS8z/OuAl2Qo4ek5u5YwmRn5iHcGpN55K7N1+1ZttQkef
rX4OdGYGpSK8RY2/970HucAuAHfyXUYrZ61eVWrH5PK7A8vPl74iwsGyabD2XlJ/iaVol6UwcCsX
vFXmhMhq18cbkcX/9KECM0jaCa+GQpcVT+Uskks0pO8jwFJIvpOXYOUuhlPjBuEJ+6K11Fc6AcRP
t8/VhcZlLbsqzfXNf9NZzFBRYAgZQJxM07XgtA5DHKt8GwfAEUYJuGxnVjt3/r8ofu3bQolf85s3
5/AbDOkXCRMirS374vC7jJVeObmB3FtpSkFxT1GxsW6BLhQrApybfu8dNMrHcw1TYKn/EJaE/VeR
W5S17hiQluX6UQ3ZyMcILalw09Px569B2nIPrqUrXNjdYHpo51JAXpx0J76uyjSzz0dHCj8h8ugg
By2ZGGsorbIKUbGp2M3zNavxO9vUaH/BblSWjp3+wKDYz5vMXW6wumDh+gahWF8/9GH41eaOqgg2
YFrAjNivvNoD4EjtxfrPJd9js8B1jrcW4P00+6KQwF4YI71GRY62B2prYHhaW3OsS/YbFTIDa+uN
jLo6qk1FvRpVRcOHwKz2J/1taIT8GdXDSN+jxmktgE1Z4K2e6PNsPX6CZMXoivcXLRO/FS+Szu9F
Vn0prOsYAwrE8jQy+ZhGY9vPnJXjmAVnLNnzvclBKNSJMSlEMdUeTTcoCVt09AzV0gGsYsrPAPz1
1gMICeRxNqX/jEICmth9+WlSUq2kXDUJRr8LmcUvK+oPlIjohkLttoR2u3sZTpt3Vst9Lvk1DpWj
X6aSNZTexKtHBMAIjcpdurQOLlfVokjKpnt+DsoXUYXB9PvGEO8oGPSQydB83KDPDN9nF+NLJVEG
8019Yzb9OIcgbbe2iSmG2HGDU/Aybo1fzDQ9q0wVUeX9r967jq2eR1zSQdlXue00tC6mPKFsGKTU
h+NuCsWDNfoKwJUriQazP6SZ0piB1Qw2u1kVsTCMDLUiGW3V7zucZ9KgRuEX3jANqV2fgPRffOjz
JT7qJX9tih0Kp1O8u/SOHijazABRUoLXwFG9W+/5wUUOtpV+PtVGKy8ShrPFtL7t1SmXw3fhNfx/
oHH1CRZJe5nOn10MKc5UW2pk5+4ehc6mEyOgPpWO6DGJRFUGICVjuVcPYHRVLOFGJuHXBBghZifW
oU7pEz7Ku32rHF3KzUty2tGfrcTOJcLQP7Mr4/RkQZvjzVlO3RyzUqPMKxFJPzA+P8t32IxLtvMB
yNso0T0r55SzvSI9bYFFoe2EwNzkEPMi9QpmkJsSjf/S2Pzloy8B2WQkN25/MONBvbHX+cs350PZ
j6nEjpzBGVX3Wt1IV3yBxGLbGqAcjkEUwYzL+YF7Y/EZ7tiEPR/hiXiiqQuE2vsZMSjQtI/7L9yZ
DCuW2AJJgwfIJz6w+R2ymGD/NplLBQ+GEbIeTNHYp7f5rAxT6u9c9D/5VQ0tlxQzrkM8PEfoc7oO
m0sPjRXXkDBOERqt+jMi2eUbi3VwejnFi46plQXjUWLR8n6dl4oW1A1BfPLqOU0hlYGl45+Pc1iR
51oU1MAD5F63KFfgZx5yM/W4w7ayfUxspXFKHln0q1qWFukYzEt7SQ2BzhToP6CHkUwYskSPQmCz
a88q/dmIJKKVRqXJOhkTAt4dyWWdvvRHZiOa39xoux+/Y0Nu6LcysACgvi6Z+pfMmwmO4hAJXHvL
6Wwp7efIqU3xD82it+pCyj18j11L8Oh9YLQbZwhN7XR7LGE4dhoHJcL+UBr6AGfjuBjJQgAfyf7F
az31HZNbkZoVYz8vpsIzkh2wscxCz6l2Nr8LUL752HHd8gjBCmpQZxDmT3ioPJ++Fykm2pe+8RYO
Kub27an8dxRyDWoJtnWXB5ExKRXNKP8moAyxn9UyZD8QWkuUDHkjFcquVsSpamRWRd3U3P6lY2Ro
ajx9DFA5lpkIuwJJHvbXueqAI1B6sW1eZG0EgzpK1RWaMo7xiTerAT1z0OaCDntilOkVhQrDbfCf
CH02TUBG9mTQHihXbA4b1ZN/3uYWT23vFqqlSaB9YsE2Icb1II5GV11nCG7hQJ8V8gidcRUejcRp
IcuB1JmQvjP+H/405Ip2wqqC5hHRnyqf0IXkyQ7LIICgVpTMw4kFbqgqjsApGsuxOPXHFo4HY5NT
18zRbC3EYJwKHb0cvRHeTJ3lvyTeX0smH31WOE+yVQuQPHYtePYZKgD7W5jq9k/tJ+6If3YAkGTx
BIvYXHRgE9YjdqXnEJYK87sGc3eoc2xaFeiZ9NDlyucJFAcsjtWUHOFKQNZbM3JyJXevhgU/F/8G
3w6b7zoVZTmzPorrOBRRWpf2id9tG4/sn46xyUreiQJhHSHGyFfaH8j8lo4OmiqBsn0UuPte6ZZc
6LvTW+peOsQBEtrO6znsdeKSWsFlrc8C8HLu7nthhbANJjDqEFMyazkbYOsJm6moCdKenKr7D9K3
Z/dmn/LN+ZCYusibQkNUbQwJhg60JHOnGYJd/2sBrs5dfXi/ec5blEzBVrpAGGy8GPo6g+cMjpur
w3qnID3NvBjXN6GhBX6FsAoQ3NbeWgcdZWiDMhPTMjhHmtEKTv6D/WJjUmKoAg1T0fddMQtnROQn
uOZ/LLamZlf4klxFVPEJ8Z3R94FuBfuEU6IZ/cW9ugezayFiUhda9r5Kf4gdCbpJi++OLGCZnxw/
jv8ZWIV1GAc7P0gaPOyRW6DKX6enApyyZ4z7FbYfOtC1AjDRcyM9Wqbxj0jGJ12P4H0bZ4Q97qlb
JoLc5nI5Ig+G4Eqh4Ftu1ytLo75uzKvXgYw6tLI0nFxmkGqtvLPNSxBkt1KaOv1OPARBU8ni57fj
O1CK/znHovNFjRD8q63T4CTpRjm6YXILZeAbIz6pUkQ0xKwpDfHn5QPU8wJvN++pXNmOmTS/tzmF
2F/XuMDnI+lk5TmU1zoQMKRG9waWS/naJFr/y9Sc8vx7LsBW+B3U+DvTNKeuoXyRvPNjFKh6gK2H
HlqEq8TYJnEFPcRA7b+S0UuyL8LgJAkOA1lgBrBCxV2kE+tQQ8wGROalct/rdXj5aqItBfnqDDpV
k4D1R5APz1/5nD04hnyGjzIMRmRPISdeE3BDknHQ3fHMynQi8RZYOEFu2Vx8bSaI5aVerotOR6+j
EDXMCyt0HTqyrUKAPhpbVHYFOJ05OUtZs23Mh2zniQP2jLWbqkaDuEXztGZVukPcx+mg78hiOMYZ
fRZTcnNSF0U3aXi6PXWwTEFsVHaQbgNik+nQ75sLdb5+31zZFGZRc2mGZPof4E2QioPbV7NV0AFQ
R/MgJDS32ajGfvFUC+1e50mn1drmqbJlhTR/Gv9XxwF3Y19n3orm3TR+Fc7N0r98d6kMauAMGdxY
N3oGtXsNra50R/gRbEbtF4ZzzEauRyg9/ZYEY4GcRo2FWBaCqybdz+C+hrY+BBsW6vbl79r9v4wl
6U3bBO/EVd349hwmY6kyTVbhxOGToGnLlieh1fcW84qsi8TzThNKkAFiRIVbwwMfSdyhFBJeBBUr
wrwFSZkHAapyruo+3yyOljb9a5eMALz7hWto0Fv/5yBBZiWBmUE5bCB40v+NQi7kPVrCUPCeo6pA
xBh/B0pCfAbvJe5j9P3yO+irDKK8LGYpYc1AYAUSJDtconb1GC3GNv4vozF57IPEEpJxsIP44Ntz
N/k3f1kzA+mSiWFxObCOkn7QGKY142DoGhyOVaN8QBGwLBIPGPmHSClH2iWnCvYb1ISM+ioGieua
YDXSMonc48DrTTQnPIqqR4TpPCiIJuDjm3w3uTb653ny/s1zPEoIIr/VZnweE3NsljHQcuXxb57s
9lis++xhugMCaxuUyle79dxN1/OLq2fkD9GchrzukUpefnI5lGrTfCqfmSjiyK9eV1kIORlYIVRp
PAc/ovUO/a++42tLtilTGyGJ2tOqmnUl/VE/IGpSZ6y3cqIEP6NOubc3dZGo7wWT6C4ulVcZwFUT
jH1u5mL0wl+OkfOHtxjjAg1lN+rWnPlTP1i7+vDnA/wp2/1R6lbOH0mjougqZwLtWNJb3JzzOhEJ
Zio5i28XppOUMchbHFbSsDoIwuhV+xwGkKoJvhxzux+TusLGOr7/SXf1PW9Vcz4nZJph46Im1lRJ
WZRqmnUHtokhPwwKVvMSFcRUjYgNj8KBEsgwu5YsZh3yHPLBgtdS0UnErYhfpmBpyLJJte6DbD2K
uBbZDPo1bblDyAFiiH++220+EB4699jH9Bz2QjT59nNymFQ6Y/C3a35E7WrFlLKOi7Y/o+PwvHLy
sTBbZhI8ynjO5njtaUm4LMUftOKpE0114PzYjBdnz50GTnSBc9BROHmZV6HH+1tchEWguIQ9fSm8
GTIzv88MiBSkq1ok20SAfmdi4+x/RXNVdFxx/TwpZtUMH0Kc3peXI9qbibboKqm6Nm3sO//b+5A5
EDy4Jt5QHcqQWnVl6XpAZ0qyHg4gzPANviUwXJzWnfDrUMex50WIewORDEOGXsVs/y0WSHCGeuYI
M8yB9w42XxEC3LV1BihD+CzY1I9WZJFYl7Fc6f6FaO9akULUDfxvL8KOhP3HoNIFnAxYgRb9PIJd
f42PDOGJzuA94Rg0T3uec0LgJdCMJyLCM9V066XTSJYH2ZPioEGkzrzp5tE8/ESDw4iffchecN2L
MZOCsGR3rg3p2KuqLU3VLdS0PjF8NaMU0LhBf7+uZyvIZYE4cbPBrgUk+9mXmXDPGL4XZMBWt67n
Y2t5mFS9i9nNDlXBwoSX/mLKMzJava0zM4nULwlmikaUamyOjig6Nu4Ge4vtjKxuD4TP18C9lXk3
DXueBnz6FCcy7ZXMJGNE8rRKlsQczpAwslsILVtoXvWkncSAINUugcaBYlv5WqSYikbw9l4y6QH+
89J+HdOJjOz/maJLcT++emGKNPrJILYJZbDZLvBhfhVYQ30awv2clnXdKBvuBua+b8LoWOiuX+qe
3H9uHSDcL5dPrrEviRmI3VtYqvER0SshQSk0BipNfe4UuqAT3qnVcCXCAlox/MeVAu+vXpLgxofr
OAoFiUKtmh72Zxi5LFXJfk40Rb66VzEZnyr4cbevwRrPb2uXZCS0yJ3EAXtBzP5f5a8vchzkmSjM
hRuvGSpb0RTCGKznEvspoEdu+Y7OQyGObL/bMDBCq+zHj1BqOpDzeMdlNWD1uuW8OIHQGhTJ/fPu
CLxhYyoLEDDVaSOdQzhHukL5GAhSBqcB0vRsLGSnBlXmQgF3G1yeczC/8GmnhpS8eTd7j0dcyyGm
JtgHLY6lGvllUA2Vkc2X6LE/69nusWwxj22z6npVykSACFcCZtmIh7djX1qFBla/Z60Cbb6yNM0w
/0FEmXUp6j2JCjN8AUmGTItbxZBKXqStgvQbmtKbCTNopYY2YT2jExC8hJH1FLDnxrQW1eiEOfWn
Tct0g0aEx1Hia9GDSZJPz8uYflNTnhkQGjbEQVCHzexYraiLIrhkS6T9co3LCXIN+pidgSU4LvOZ
n/DKMm2E7UJ0ddc0gBpfl6r3rwrsT8hvgw6WbXpIQIfn4pk7AUrtT8kFZZkCr3nEh3kYm8BnErF5
3274xqrdip/CHuuJG6x/obyFuCSWukO0lU84pyF3Vc//ga+Al7wmFCoH38gVxZFWPE11FLVtXM+Y
e5IkMAubWbNKfip5D9cu5VJh+KNIjsI4rbRuM6C+W7SYBw841b3rLswSOW3Wq+gRVodRv2rWU1kW
daluqSZXo2oxRvujk2QCx1zgj7ukV7mS1+hETsqtaxM/2Dl08WwhKIS84tyvqYvN5SI+sqIM1GET
YzrzLKxEKztlrbZRKnAfR2L7ZliRB/n7XZAQv1L7ocCKoT8lxz6AjncfDBD3Bpaa5ExGQ6QWtAaC
heKKROfPiI6j6JjfkM+QonrQ9uxOlNvkoxdwC5iMHf67jYm0GA7BYTsXQWY0D/0DZZNB7pEnFnrZ
GF2MSAYeuWIf9tIZVVP7QjjsrED5Z4L3rv71942OdxbRxVqflBuQCva7rekTLnz5FP/VLj5SvTOA
GzOaanKF5IAxP2+ITSCA68oI+Q7Rkkm6CEMXnzbF8vEk9AwqzOXZQgbH+cHXnUkPKktt4jUFoSmJ
HPnILdq7YNTfucXKTXOvS6Aox1U/RcVP69CIIBz6yEU6BFjQuUBZj27Iyp0fBC/H0Mr1jEA5ONeg
6y/NMzveN5u2rHSMrJnNieWUfticUr1/+H7wKBa5No4Xk6m8Ay24vNl4603rTCpzxfqCFgZ3O+7m
d+KmYJi1s5+cHrTd6FT3vaY7gsQOPUY/Yz4jqHxwq5gGKNSg7aaXCqmaWqrt2yfQgmG2L7Eqs0Po
l6F/X8TKYKAe7afaMdedFzK0wGdoivFoHKZyNQNIAwKSdd2C0/SWMVOcF/T2BIC0nDscNwo/5t/+
TGKy0Frbit9k7DIu/sg4GGwK+lIbEVXNSJ1XT1xwV6p14z6Y1tNBAbmaeiZmfGE3r5Fxq6WVIkqe
WzvkxjN2oqbKqFWs86FKDaxqtscnx4VBXa9q1F/i0mAF7kn7rM0xuTCZaRefg8qxfhcrJrPdum1S
V33Qkb26Q34vrl44b07NUCwK1WVmjJ5kCO6uCO7Duz9Urn7H0fL9/vDBomftEkSLhIAZ6TZWnvxr
teAyV/8K+Ki56JIgFssr2MvwQm/koUX3ZSvA/7Q5QqXDo9+uScij2FNjuv3mfgAhPhBiVDtG4/Hv
nSl523YHgO4Y8aRZ2tcTFE9bPfdiWVppJD04uO3l3PYcU8duhe8jokn/LoPtndpeTrWkh10Wx81R
mo5sxLO98s4W3B4RY4P7IVF7pufRH7BwuPE7oJpE8l/hYKYeDydfJ+2pPBT4YXAayw0ItxZujvJe
AiGKY5ABvu6bnRLy2h+CSpna8gM6GCkwrF8xTPP3GtgYifwW2q772trvyDCGGQMXK4KAQxQiW/lx
1TmIGOuMOg66Dg6U0iGqq6TQPF7Tdy2AVJlqP7ydwoZrMrgKNoHLAh6JBUWaxOA1IGWzpOdWNd3H
VePziHkO/n8YxhgO1duLVEknLJHqMDtpznwldZXH0xqsYMrIEa5LBb0G4kJbuqZcJcVp/kKYryXa
2mN5pB33Pn0ZQee8hiHbv2d/lhuiSpY1H4vNJs2PZbMft76/1nUIMfffpDlbu7+oD/ShIAoifeog
I9f1TC6QkzyEGvV7GuTDVoEjc9rbisllyBKJ6yAqHu4/d8FcaVIXBgDbXmT0sFpi+XED9TISrajM
7WMAOczR+d0cLzNO5m+tEPZXEYFm+bRnSG7W7pxGuNwkT1ulzRo/hefkVjNi0MYEYQfgvbTLr+xG
KZQPUitV/x+rKekPflSJFoXDhH83qopnzENiNfHCfhRE5Rm+kLxp3stcKrLJKLmbLDDKrhX0mnb6
aG/AKF1SQrF5wNvxYer7IXVaV1OagBbZdiUxgW7Jv5uoRyL0YdNUZl7FzIVxIMBy2UmHuE/1Hwr7
D5z7lzcMCuwp390UNi8XuDoWqrn0kSAkUz71CHFelvUx6ldSBencTbZNVKxKFQ4hGPuUySI2I8IV
lhCqOFcDy5InH5ngp6XHHFPDRnqZQzGsyb6hHM4hZK+ixcux0RSwwFpdUODLBxyx2S7LXxTKh/BU
9ORz7E3574kkY2L4iyeeOHgw8ETGIGu2T5GGTtMZJ3848zh5Eh+Z65PObtakS6rsumDGuJX+vBzU
2/zkrGKZdsJx3zUrOdXTbOMEQAnS6Cuiv0pbPJTnaHOrEmi6q72t+4+ElEd+y9JDBUP5AdV91Xde
kadq1Bl512tzsQc0+TRj6EvSUUWxPbEEZEtcGkuvik5xo7L3kSHHCBw0ydfj0fhcmrOIEj3F0PBB
qcrbDKoL2meTCM1ka7mTX2k4xIcxxaDzGi2qsZBPxBIXjA1qLtAFNMB0Ost70I27pYwJPS1EOhBF
6QbetzMxkcGqhkVwqpFHq9skGYN/C9d+UiRpjN4p5a/jdY5eTTYQRktKMygQpTa0CZKfoipLdnr0
FFa3pQaXijFyB6Zzajhd4sBoJJoKQIVkx4OkRIqrYIrUPeb2SsFS0+zm32vQ8q0M5LJsRwhgVMiv
U+9ru2oSuo0FBh7SgOxPQL1CXARH+rW2/TfxiXB0xZCDV5M8dDyp4uM1tVMgObRKq9tYB1LKB4v+
dCw9WHDsr43lyKBLD0WhvD9dkCy3b824ZSbj3j1qkLGC73iKyUqZBKxes61o8Hw02z1/+0zF9FC6
fRXDwa3eEZiBkAZXj8TFOuS1HIcA+W/UZal1UZgzZDiRxhobrUfDFXczuhWDGMgk9qrZ/Rk3QYWQ
LZpoBRGQosBTsvl5eXNbsLRqk7t5VHkclKxAQtjQ6Y4So8ohUxAzuIWcC+wYJTvv+5o+saMrlBAH
upyUghHxLIDadCjLnrzayDQN8YoPwIzh0FPfmdS/k+ppLJc9kveXfB4pKN8aPxTok67cChnTGoFH
jaGVrmLTJDBHiPRKq0ENe1SJruY4h5ntqI3Q54cAwKGFFrLSMhngkIPaefbgjuXKeU/d3Mxz3UTh
RPWNoOKonV7lbRrBsF7RLKjqrrzQshMJw6rI/YmZekLB7COsc21LvzjbaaXKvNah1I2n9A3FmKSU
dWcbiy+Q14tVIrUzkjUTXmUeZ1FS43QWQPl9F3SVU8cr4iHO6zgL6T46g3mHWeq3bOx3ZUbf93tn
yTYLQ6ZCrEpzWaDEErbF20bnoCMnz3V0aXJ7ZCTcyP41smXyPHvAwBp/w2gVn24CZi9IwQVkJQBc
qNOnGZSovq15n2STcr+ZzZ5MEw0155trufh89+VvoAXtOSs9gkkjZXGI2wlPknOOfqOsjyf6Ps/0
mt+zAuScrEZDsmL2ABdpc9s9LiqcQelusSNwz5CyLv45EgQfi/HvTsHCkxp4pWfwCxPsFlSa+OF+
/iCcfqm0MNfPIMoAwDJs6lSYz1S1V0RWhlyCS96eYSi2BAbDQAup2q+cu/TbtQP93N55JfMiFWIG
H0+9DsvpMfGIhMkkXs87Vy7rjqHlKyl9e/jxrboqhHKvQwgyP+OgW7N6llVOOb3tgf0LqgH1VwZj
LzYIGEeWEZsuT5PUYBnBF17+JpiAOuCnlVHAodtj7e/p7p0Xp2WzZ09DtU2tk4aqMF0doGeDR8SH
fNwV9KX8OxiHlVHruDMjax3Ib3Hf9WSIYq6+Wqdb32v53JEXOzbxR6WHRidwcYoZAjZiUT+q8Mhp
FH9i218TgKMpgxJhhPpKf0XtJI+qY4lI6mY3SdymEN0wTBgNePNvGHuTD6jETFkxlMw0xU02a7BW
u56td3/ehSbONIZrpkzyCwQPG+7jNN27LhSik4TNMcojpCOGvjCQnSw8q6RP3V9NVS0hPlny/CEY
rwJjGcCpfQZKCPxqMWUTV0mzHNz7m1Q+Ua59f/F7uYXUXkwWJ+jKvUEWUnMhgooFuEI8O9LQZnXD
M1fMce4x6sloZg+NN5gq0rzQXUTYSDiUOyFKsuMKtOcZxiZWQBk1cdPBbW1BSEHulVziCboOjTAa
u4OQJjS3IjmkbDDRKifcP5VvlCgXTi1jInR1fLknMuEYEqztRD1qzb421ppqEoG4zY5YdFzPorW7
8Ejr5g7wtb2dEMAyZ1JASx+6dSaOw63zGeO4rdGSu9ZAq6KPjSM8dusJcVdHWeaynW2Ikm9h55fC
OR2XvdpR+7KgiZBr8h7hXdyKVPeiuC5tWOxC6/O3Hr9IdzVia+E+OEwlslwc16W3kliYQcYZAHue
XeXNVXNZ9NxGFWgheLCCYwIxi7X6CwOyibPm6ulojt5ClQgtVQX6oLa6J9Trhvok48puUsmLc/JD
/DDpzafv7gCEQ44+eQh7jBfpdWIIh4EsEAGhM5s8KZO8aDKUABLCU2LzmfjORBBhhDj+UOo8+ECL
toroYxlrp9AF3SqM4WdFtHZBd5t9WpYzjaqEOBeq0/Ue0Rngjy5paVq+WsiCnLqc/J3v10Hcp+a5
0yuk1hfjPBJ3s6WzKCIYZWY+fjbq9QRCktI01gY5vw1jO5q3Edq+sKk+3prnVecZhg4VKX/D4LLu
Y/YUI+jVj+QOXv74RRhJE9/CCMSUBVtjyueBJ8EpgoeXd9t+sEeEfmnFXQN/TLkr1BDptAkHUr+A
O/U1dIXWgFBQJTlkzHXgjBhb+lIZXenvSyDCp7a/jgIn0Jn0e/UVn9C0fMxl1ekECHI28oa8R/7f
LmuwEpH7TJRrQLIrD3j8yptmufAhos/UCFgyFX8rPCIJoNGpp+VPIBinbHVsmLVvmoFbL6DS+ezM
NOOS5wW9NC1nHej2VjTECYDak4IErKL549aHV5ukkOmhQOnbybqF0tB5SETa279hiEyh3XWAOTyi
zc+WWfahsbjr4JZo0HiIsbHWxit2iLwZP4lEfl4E+YWi9PWQHtYRtQ0iF3+1KgeNiZ7MgbvpnTWl
RIqJ/UQOAdnnwzDbf+24kpXj5inrS2gsj0HFtsCMuqZbgEzQal2E6tNduf9p7dhcbp/zW5CuEAl7
8++DF1w97PNocsosCU5DWhKrFJKBu42ucg1Dh14eg7gJG7FhHY2SE36tlWj9cDPzzygeTqUlk3fO
h9now1NZE59rqdDDEiEog0dAkA2hEXVisvc2LB8i0E9dBQcdbziaU1/fSajZwr2Quy+WowtjoLSk
/KATpK+UgvhwUcj+cddJnDNYZ5Gpp5mVA0Hsac409StpwEC08K+vHwtEvyzo4YvMRVkPs8qvSoV3
1yoMEIB4WweRWtFSQSv7lGX61wuDR7zOU5vfGuWNZvUwoShkh1VflszJ5hxEguIkKnZb8TN4+TUi
oJPyDBCGSkNjWlrPZqUAejPuj+TrIbeYRfroKRVegyf7xjVZf3B0SEXZkbfOilvWjYIhowQafkp9
/yGOtt86g+2Tolf4rSqQEGf7HuLn3EJtDHL0O8kzcow6/8JRfXEXToTJqtDHgvFQ9Ddtae5TI8W4
tiByBmNwevy3FLAIn2kvwZk+g2tJ9k80bIWIpJwm7nJEBo1hKi+lRewP6iEefM8wUyQh0u3zsPz/
lNK6y+OpgdSl0s4BMnEBsuIcqjvBFrc2yfijz4NcVKOyNXICJ7KoVz0P8YbjktbFSFUCmkT2EoYE
AdnPbxAyjrauLfENBTaFFY9iV77gSHLs+wf3DQd68ri6tPfkB+SBNHAfs6DTEv83IIzMaUDuWjUL
B0hhdCbj9/9lJleL6zfPSshuSwjROMiGUZ6PIm6KAzRhunbdYkAEVE6FxNmVHzKt6V3ymngSiGR8
6HJpjqp7MVnwWvQoAher3aBedUsNTraYqA+r4Lce9ds4DSfHIfixjn7wJJjPZQu0X1SXG5BfvJOf
kNXYdCYQE6KzFRAb1H/ck7KMYDq9hAeWeREtMsjsYYLQfBWNZvWXzHIn0YDf3AMVGkRrli5/W8Qq
I8aRd4Hf6E6B9zkbLU4nt6OhNXcW1UX/VErLPrHQNYzx0MS8kM4bknRrZ0hCUvuJo1DnaO3BcAa0
YceWIcU5hYQs5oSEPCzwOTOOVFSrmk2ifB8DCMw38NWn/HS3CQukAIEH98pcUqy5nG3foUXVE5qy
V85JX1dt3ZDM/V4NtGCrqNGNRzXHBO4W9Db/sSJwUP94w47RWnMvNUMZXoS49rA9Tc7MLdReJDxx
DtajtHSftWSgn9jvZjk2zJNwz4kaf30yavT7r7+Ql2LuA8WKGa0dzbGc3tCIhww/UcTH+2hOFe4t
McDIFsxU8gr3mHArHj+wHL/LWPhTD43U8T5/BJ4p0i3A49sIvX2Vj/wbwOacFok6AclekoFMHJKc
yU2LXn0hzwcWXNm3nD9Aju3OXfPjSQlLBcYftJGa2Z7hY6+pohPDmWhwnHNP4uQ0cn8JTxIZHFm7
jnFpdFbJ09lVOfwcliK8WubIbR02yRqfSLkgZUv5QIowbhqk9Otcd+iVyNQhh9lPvM2VouuPqb2v
8PhTpD4ETKF3muIMIwO5BPigmDSGWroNxc74Zuz917DuFn4mKr6+0XeUNAmHf3fLOVtxBSV0kOhD
4nqrh5c2YlKXuKlk5f6j0lp7uf1znahfG0QfhVE3QAUl0OLUj3/h0J9FRaOlxWy/k4tjbLlB4ecC
bbdne7vzK5fLDdc40NLT2CJyOYhbsDJ7ECHsMrSMc23Faw2SWMP8FXge+nFczEC9xmGauKhEpzKc
IPxgXnrlmr/HV9aesC0ECyQKa3dmb9cZHZftsM9Og+C46+ErMtrKI6ivm9t5QomEJGs0hfv7JQpd
rhrcfQ6JjJ+zCnUwW+ygFnoohmG36pmJH84eRd6Ck5G1mLNNKvbFgj0YKDX4ePhusx+BOj1gPeyc
dTbPh1oE25wwhx2cM6lAsHwzGwM6Pu2BLAWpX0IPn9VG+DcreMKREge38XCmbFu/2RK0FYmZdljv
XeL88ga8YiAR1OOGyZ7W2EyrW2rjrgO93Tev1am/K43pys0a+LDYwGkOIdb+fWe97/iKB2SB8CzK
++Qte9b9gf2f6vxx4OsdcdLrBeQI0um1CFHKoE8cJwP9/XCc7QzviFfaFeuiyGmzAfsWTuoS6uj6
/XafywxBSxLKYTterC2pZBBXtoH29OujksKAe5NRfj+og4r5ljTLMUuAPmIJ0VI/r2NbvgtZVwkg
azZ0WusKUprYxMn9ZsZsm/S6vJwK8Orlypv6Hk/SU41SAxgHaYp8i1RMyEACackmmHUS5BPoEZEM
zvGsTyTN2yZqicci4no9DZj7kCE15uEnHntemC7Gl2pjM3d1MGiGMxc/ZG1eDZXgjQKEyJDXYrv5
Wyf6kLuEIbS2EiGO+zSYDMYkwVBgAMhkIHl6Ex77/ybFOxt071bXUXtdkVyWMvtBPdemAF/iN5OX
ZtQ9fbs8vlHRXAm7Wd/mKfygUfGk5XI26Pf1PD+lIwQ9ZOfx8Nk4nf3L1YZrhw8Gp4h0H1G+OZlt
TD+f05uYW6zVZ8g+ZPcIYmv8RntLJpTBdme19a5cHDk8DEwVhEIdyXDRdl9s2U/WP5tklUTqlX/X
3EmQF3O6h/Op0ctuI6egzFPGFPnt6aIMza899fzP1WmYGS85dkKQy+iTapf2tDsLI8x+GEIdmq/Z
1MLLkXK5kvikFBoKLqSLyd/Wcgror8cA8zOnlz3rPIOA1P2NrcvH6/gqZ70AHs98r4b/0z2+6yXA
qC3aVUoU20VLbsciQbuP5J/pgkh9F8FMc5f8qK8jfgv4bhwdahWK8dSiYRwq18tVfQPXfmPt0KeN
uOfvJR5h+UNnjmp/nVcFmu7TZNc3nDXL0zkgm17buQ3EHobza0p0Z8nAA9/FsxWgmceTtaT3uCWl
1DwtgP2gg8x0I4PtYfvD4a+E9j4a4zxrYKpymvAnkzCcwsxD3EGow/ZNeAGZuwMbcDlUSyOcoLtp
X6X14QlNIf1gr42ND1MYfWy3ag7RbYzFyWCjgHTHa7/rDt4YhfVu3oXxw9BfS8wtFpbpYJvz66Qb
li46URsT0OWDBbjlGK72xj/BHzseHh6CZ4M2592ndCKVWHzHzgmJSOszZddmqFmvj5CDZ1wgdwUE
76CenSGqKLxVyhpV6F7jh1ZkGKsPZTkdVhOSvGOOx0Wane3IcygOuM56nFTnG52oP47WNf1VwfEw
ah12PqC2ZlI1b9mJjAeafkrYZH6OCcFNOgpSXnrmon4Efsfa2+P58u8RH8+H72SvKmYNBpKlDVXj
OADHNvOajtYX/mn71CaCsQAaTGVVIYZ6NxUn/78PwRKf34omTeoQj5i3haSJPEVSCkrR3mySRcCo
wL/mj0br3HVcaa54opntNQSuoq8a2NHypfWk8nbTj9fJg7RP1vFJCaCP/6CaV9Z886nqeaAsHT4A
FJKiAlrrHmPXi5qdmDBgoBrh9KZoNDLOPXDJx3HMkte0Wg9+CKnIk2lABx01KIKcBbrfI1Ab5NR2
2CbIm2Jz3NIgSLGlGzS4dNq1m61GXS6EAjKQGw4Xh8Wyy+7QsJY8VZK3S05339jatQSSzc5Dj9Ca
GN+DElo3GE0YIJqzx0YBpuYCGIvoncMQ4W9ce4KdjA2f5XTKLpSBV8mZObh3gAd9AUL3kHXi7Ca9
fyir+O9LhZ4QKIhmNQ51U4R27xRGnqqd4eZ3RpJab9uMJul78E4RDE+UbV834MJwClEuZRc/II6Z
OXTQ8+HYXvHB+lzGCT6j6eGn5AKgNgRgP8bj91DtgpMeLRCUNwg/KXdY3Zx0W/516DcZ/j70cXBc
BSz4sdyNnS9F9o2N8l6ZSGlvzDwlgeg7FTP/ltznf6UUqY0bWvPdgCjN35PwlLW26Cr20UR29rQV
WKdKUnPOE8FiQoi6CK3+RbxiG36WmUc2PDA8geoblNevoLCGfTswTJ93ruZebysUBF3dMGnWfd07
BC4DxTmBhNOiEo7wl8X449X66mInOh6tEMmQd2qsSzeC+IxAMUUFb80hbY3nVt/+QfYCPr+f4EIR
kagLIBkgKuWaYsnySCH5tQPip44JaJqsRPNVFBsOHw8/GfybzKSWWH3FIMroStYik9nG+C4ElkUd
spFk7i0vkFX/SYMNNIYpBG9oIJUwmMAqD+8jcTvxXiwgHxrQNLxmXpziB0tNPJZheZ4N94Np/wjc
ZciYFSlceu+Mt3tGMJ/704Tty2cL/b3FFvzHGINttLCIvLeDkDV4Ldo0HEmWqDZbZrq44MNc3TEi
4pwGnPbejtCywpfVEd327AYYF5PIjgwXu/MFLwX2EDqrsrKeP9byvloEQp7g4qmttRnbVQqAg7p5
EwmdPTnou9db3/3L05pOmXp6GDy6MhH2O2WrDRRWoWJ+h1mkLmbxHlxM+9jftrD59dLUcKSsQxLF
ceAzamstr7PjO2ujNZIYOAadBlB/7SLW9RKqHOpY8mDfYWFWKCxYEgIpvUcpz28tDL2GapdlRYDO
kOrpxfa4j868J7nwmmPgDFZb08xE+fcX3yy2JtTTTDgRXDo1J/qLAMJICkBss0cCwcf5Kn05tYLt
bMTdcUdkH18uJxTcDi13mzv0dbR30CbRlMMPIcd1xzhsqWZYjEdEqnRwydoilfRs7+Vw6dDEQXZB
VmI6wuTmz5xiPnh9R31c+31LtEjVZteas7r+NPOcbxIhFTAENN8xkUF0DDd5iovmrhg3XuHHdN4S
G2/DEnfwRTOlAKOP95h7uNerp2pr9n8clzhTdXgBA+eQUwP9lspz0K63tCjfkU8yUiS1RsgpFXdQ
OXQV8Nmy/XqaKVH542gOSlcFWC9WU6PEzHqXVffotvC5A5DoBvyag+liybHDslOq9XR4r7X81EKQ
W0pWFakcBc7r95fWqxqn9utqKrvzZ8twMx9xfxq9ZI1XthIjI1W1rwioetbTEJyJnvDZXRXpmqE6
vdmjQK/s2KStqJWErak84RHlC3r1KGca6afVI9hqIyC+A7R2PNvGH8fLHfQ2nbHMJ6ZgK7iLFaOq
zPqjbD48ojy6CRnuUIsJ2fXK+RRn47CQwfSlyoN4v/rZx10Re0ZDmdGppe1xJkN1TXRT6NVnpsoZ
inRXjfWMzEQNhfdsZr0CvO1mnVDZrBlzKXo8uiAkja+kbTwbOIS8BjZo4H8KaT3+rMAkHLPyNMOB
R47amhmYe2OsCgzJJ/i1pXi5FPV4Hn7XJ9uy0JMNQ8G5ytPLq8WxjFpA8axnrTfzXdc7ceM8xHlB
Ginebw3lbS3dNUxBL3MO8pLc3Fj8mjTOT8hK5A0I8N1lCag1vO/cJYN1tFkGcp6gii3RChihCA2u
n57vNWEr0QKghImsD0Im/iRu+EI/lNY3djJDY7E4Aq2W+VaTS5qta70fceW9KP3Jvh50Q0bnL+tl
4Z+jGzl0IWtcwn5EZ58JVau8Q5RzSelD8g+lQjw0U0/BG4Ex0rj3TWh2RVIvnEQTef7g9QsHqJEv
d9T5aASl0NxI+zSgDT6vpqRfJLtzy3pw5u4bsKw2bU0pZVdVniO0imUMfQ6q2mpyyWTAtDhrNdEm
H7LJt8bP2VFtSgHpzuowqmInLQJcqnKeKfztcTGtZmXsDbGav0BxxckS9LjgeJffRYZRb9kXbHok
peg+C5vuKKZY4BEevxWduY2v13+Ny+RxoQnfGKWGNiOuSOyisbD3B9z7gPVRJ4tYHILUedSYMIUW
0eTKMSYyf76TiXK9ZtH5WvugCMKIbRQYMwX0hPeOOmz6hPr02C3p7zzNIQ6w0p8GzbpG1Zt8jWb1
yrcWwaXF/lb78/L0d0Oo3gt9Rl9aCbaER1SR2CM9kr/hDukO6KiB/8vWpQHTydZNOdhKsVqq4apq
B9QkCzGwiAbDsAw4uDqVSzi6WJoSqMjyCXyLlWL6ji8wTOJO1HsNDjI5bF1uaa0GupWzdd3tBmIB
JnaDpnuITna/zXBc2YYlMD5yIdgNB3Yjxzp8D377UirgUAOdZtX6THxt1H1Htt47edGPBrQ6my61
Lba13nfrw7qSIz3nPLMvaUJvITxo3ueEQuwB7Mv7A2+T2s5miiC5i5Oi45w255tRDKzwbPgqUN4I
GpeioGA6F1bVuDvFqIuriU+5ISpEpv95FsyUb3L9JcTq5PwhCBTdtnpgEo51sZkAC2Km/htcM3lN
1gMOIQkAQQdklM0ztnYcEsLHcyDRN3hEZ8rqN4xeX4aaNgcWPnzosHpoZnEFaGpxVfP0l0m9NUZT
Ab3+wwPJKQgLQj/8cD7QXU5uJQVZZ1tXwKR2Mf2fvxrmzOQbZuT28NT7nX3GjtjPew3GWJuNtnXc
wo/rIRJm3cf1i8r/7XeCXpsjOwBigIQtHwxfyi/p1BgzKE4Uc7oUxw/6GGIHYvxyj3VMFDhtxo0Z
P3oM7zmONU7r98i734YwdmrFJh0uS5pICpmXeNVsmuGjjrPWnmfXFgcsVP7PtzVU9ZaXLOX+gAhu
QmmyJF28bhU5K0EHb8RSwrCPuoL7OsdKgpJ+lvoKUIxnWXwiDUik0Y+bImH5cmnadp3bBUgYoQkK
NxGzV4YvRaaqMlyXfEWg2mqDLg+J49DuQcCVjkKCJ6dOE5md+Sc6iSuLCOQrfseBlb5VLdjBTBtL
ennsktOX+/UKeXQpI2MCnovzmPyjzsN6dcB8sJ4zraQxs59t/juOxXt20jRl9HQVyqVaMR3jhKDO
7bhP3dRVMYhUsRn9FdSeWqkyknBt39lNQZ7f+7FuB8NksLsATIJRP3ArSExLqG+OVMvbuZfWbilW
7dpIxjfwMUxB0wUHCgv+V8OBRF//7I2y31QLWnF1QBjWyB+rdhpnHz1gTfcA0raChQWxwbGcvvlF
uK6VS/8aUHRS/YgTLf/BmF0NFKyPWOChvLz8SdwYk1QnBvaZTF+h1y8d2Q7oF3eQsTRyvYP198pS
kdm6DCiNi52jR+AFtxb0h1lE3tHCuokk20Qgk8ylB2wTb6JllUT5gr/KbvEMmsr6u2Lk4urW+orq
tEd65Z18CpNVewmZQm0E7jTZQ0DtiPrOB8sHtswIKfaJ6fNUz+IkveaCvMwZ4zdO7XobIdXUyyg+
Ze8Z90P3oZdE5ZMkZY4zSgqwlJfdaiWHN20C8P2HE3qWSo1J4D/sigxdEyGHYudPsYjCrg3t6iIl
CEKvdIDVlogbVEDXq2Go81D4aNmuZ5pWF7gOb29pDV1kxSA0TUPGiWNiIUMGQ9BMn9Xc9ijd8pL3
Lb4vG5ethK3LDbkRSDgQS3GM8DkpnGa2gejE+usgCMgnCwKvGrt2g8B1I/wN3ErCyT3AHwD6IKVG
W3n/NVV2qpxBUqsD/57a89s4U7WwDPwlOkNA10c1tp+DbGzlMUMsOm1F7eTzP1oGs0E5TR3aIrt3
xmB2teBqE11OeMXrOfwydDxwXgrc0zjGysHiFAmbLej9MXuMmvbhuF/+pf01VB3ym6TEOjGwpPTf
OvGs0y9qyzDbVvaS+Iq8KzDGDmVlJci10x8772/7qM1yX1fcETlilVCcmwt0yVeuCcO3j7LWUUZW
kMZqWTly9l6a/syL6u4ssHPJgXlILw8o3qvVG0z+JV9jKJ2Voo8C4ne94qIqpDp2upvVM/Si8PXY
wRU30ZhIjWM/FLZYFf+S7uB4I2I9e/ZhUSAVfyn4IjLAxxhfJogPe9UuFMEdWBoQuoQQEvhqtONo
TJery1HoMATt+cVdUJcWuPImQaPOR6yuEOS7zAqDB0AJgBc1ff9x5u5IyurpVK5ej0OC5KuxfQUG
JINYvGLJqfcW86RlIOPw7D3A2Ny37JKTEPNvYGYch43u04T5XVZ3L2QRyAyKt0QYOkAoTvRtvaUw
d3O7avaKvEJMZLG7KxADhV/H7X+zUJYYrAclPi4mXolHlu58nSzJoWv9SwRgleTNsSvQluqNkZwA
xJ7Aa6OCTcAfC99hc/eiSYrOYPUq8sxeOLz5HY3BPeVDZi9NszfAeyqSNZQCTn18454vo9TKqZ16
Y4rmoGTOR91owlDudPmkkGBSyuPdM0pdGNZxhvg2ddgjPNarbIlJvk7DQ6SlBOpnVL3gdDdbSgXH
yj/3t41FgcX+9WJv8urlbaQLrVzplz5+tGS5Y5NpFlyhKlFO7nHyKWNtSCFGkfzxvG4AyDmcfQPJ
reN8Ag61Br3/oeQjrizGTRaPIctgpcEUW08qDqiTelHHfJg9Ms6W50S+vnEA4NVpzkfow2XMGFJX
SLsMyi92b1DWw1uvdmkGTY1gHMZwh27LUvNmpTZg9jBUiNuF8SekuyKJqbTvLIfYBJXTPV6GZXLl
BdIo3SlG6LRjf55bRJ9+vQLZON2GrmnKbxdMqXh3HDZzL8ovy3EI/ND3ViOpyoU7zjcMPLZ9X99Q
TOSKWI22Ph0kAj4k00jdgSsW40c+0qP+qYdYFBTQ5Svc56eT06JvK/6tiA4MixTERCnXnf7ps5iE
ZKI2ig40TtWXYlxSz1TW7AGLDaDqa6rWSyhnKBT4fZg21EijyeZfmlekMSpJb+Ercj4dMSuyXzMN
9nEE81ObNQRmz7vKEVELkAxayfGpyiuuwTxIDam0gahrxu3kKeq9wlMgn8k5moe58yvDyHj6Jy4a
PptISxBgfMbZn78t8N0dwoNLtzdisecUX/ib7vTP8YSSwYm2BfObIfGWNywkJxOgRzRuYdXDmmds
dmVxLK3J7JL6vAhd+UzjhOQU1YzeQZ9T2GNifN6ew+8SLmDv2q+139MrJB3YOYCDwpYlqqoMnE86
+Bq/GQVabVMyfl2EIhmrHVNv+1wBcrLfpm6GmD2nMfmTlkd3rFSr2MeLoF5IjOks9kdJomRDtjqD
wfk6pNREEj03h4jfQO601Yq0x0JZ/gfY9qE8g9vIuAo48ylIBZLJIIzxLl9Km9XeTjlJ6NW3eZtp
j7ebMG3Z8Utj1CTWx9+jviHy+WgMalhAQm3bSSgI6oPxBfxRwbqRN3KqH/HLGXaQO465CdrF2ixN
UEpJpSIK6511BNllwznOLr7lAu/5YXr5Mhcj1G53qN7JVUJ+/10h8SE5UEBXnFAFqEcmVNGxFnvj
90jJbJ02QW/1AHfVVcS0lBIjirIM42Yuw9QdnUQ73YQpjoroc88nAiuSGs9kOUqObKpg6k/FoTm6
bb++hQdyxQ1ojPs8AlHWGKi0GaI7jd9UyiqF+J+YYlMgglAZpa6C43VmKijHsyJHjXypheTrb6mc
suGT27dvn8WnlXGqDmywRANahvd6S8un21/44rluia5ss7YMDmuZKcIAiEAzwEQOMGQGVcBVOWTx
pWBO0AMe/nUmorFaO/4TmqiIc5ehMubw2CeIne08YorqAGBxh80aO1e0xW7vJ6vd1wE4jqx9b2Lx
m2U4bjyUKLdLCK2lkJYZKOxmtNA0XYZdUvVGd17tD8p2uVqfj9GqjyG4y/sccPjsuXa+FfaD3IOo
5SYgNIYBBJ5l+UjXDXJzXyazk808v3WGysbV6djxfTzb+WNAIiuZEQn4wXbTxMCR+ixqTLfRNIx9
5jd8nva5DvtrFTLUx8FYfb4eZ3eoCfUcWPBhjwwXoj391S0F7wLKgPUxkJWWz9WmmsWFewit3JuC
LSPt19yHNFC1w9nYpppTkz5GFRjxxZSKE/pIizJJ4XZ/3ZwJToY/E4Y2EloxNso0rDRakq3Pc1W4
D5ADmIs3BynSdwHru4C2lEzoW1LywPiESp2rLPYd3Pj0WCeC4SFz+c6Jqv9jRt/ghJ7OsgnICMsM
RSHpX+igwTHRBw+NRfq9ulX1Y/AsedUXsX3Z+0lv/0qVAKiXnnIGTD9KWDSck8TMrx81b1mphY1Q
PYUGd4lJbEjadbdt6ICZpuA/qPTTAPGcP7edi0Jtn0xNP8/LMmUt8aYviuUBdJxiFJ/qK1VzS0V9
hgwdooZT7g5nuxJ0g6cDF5u1jofRGozs0wUo9ESeOZV0uzGMbW/PLjJRxHX8FkeN4exuOLIWb5u+
DiIFJxwC9ivO2s9fB0Ih6K7hRqYX/jmJiNMeyGzPqQH/a0HDXPi643QKNjbu60sTVPU04VawUX+K
Y2bNgr9/fPIsypkj+kmGW1p2XKuTI/16lryAsJrb4Ef0GuW/QQhS1GyJPw2jTWIjDnzb696csQr7
BiGJ/xQUjMP3DqHMRBtpeuBIoChNz+A3SIyqTvHOhnGcbLvuCAus8CubOtJEW7br6LSGlUq5RDH4
60/PwzjkA0u1VSnIU4RLl9yYmc08rsPpAcqL6pjCRE7ErUk7NdyZW7yw+92OM1OfLo6p0fMiKB+V
gMfwY7NajSYfrKkGNclkr/dR/9dXQLlkRp4Xics9+Xl0TjhIkt4YFXZOm7UVLcRr2mBuVixfuN2t
pUFN3KVDSVqrZTJhV2pNOmZRxmkxDeTs0/dwyg19PWtn5Ejfqp7Vd7SobiHsXyXIYAIWu1gNzGCM
gHCT3hJMRSbDRajvCY0WXcy6TvMqrjnZsgDsV8hfmX0+yDF5GQ/BBGKL+7xE/N/Z5pjGpTOek5FI
K0RMllBcyK8DMVvtjNElY775/ki6kil3EvAiaGhXyhdazWtewWQg8NTVJeQS2c7ri9oRMnaauDEF
L0DaBAJL1AgPHQ/jbONxDMDspyx1j8mKNdbTDYxhNeYH/sOlb/MAHfv+05krTKI72aFc4zgqWXV7
PTJLO31kAVbhVSNsjypl/vjk+9Jexm/Msdp+VPi0BoUprfSIJNKpQR8VE4yKDpczk877oRwy1aF5
bb5bQAkwlwHK2T/ihGZ2OJ+/oDWN3ZWTdhxcYBt0REx8HCI0JTOFaf9tUMxAMehQyNlWbquRZE/3
hKdCfSPQP1LYNNyqK2RDGTLNIsf+MZpm17T9gykHWAb6RcQyqdmda4jG3/GHIZ7XSUVV83D0smo5
2kD6qWnIvNUVUN5AaIko6rBqN2jrQOZ45VS3jV6m8vX4P2OUGE1cue+ICyGttpzNjP4E6NTzklah
ko9n3daA7ryGyJzG8n7FUssyqe39wHl8jA/WaZ77kJcYFW3BPOqxkGUv3QBEvoqY4IZU93p6tJ6l
PhVPoANZkNStS1Iv9Buo2gkPlzBI1m17ludLklnp+vYkalq+/ujmMnoooDjDV5NF1VVtYsDItc0D
xf3EOWaCzzjHBDPYe/BeQRLfAgPj9t6iETvWc3qNODWXOX4m25OrpRcvAo//2A+tsdtZ9OfMf4ls
CENqPVTIad3ScKMLGkYZ2jLW65cQd9KTuUfQzBMmyoU0+XPmzPUg4OgvPwjg02pwnbVK9rFzxdN9
TSeWGDsSmWknOtCyPeAR7hKPF3ZLDBJsBe0N21Tg0CrzIqA2QiXfanQc5+Ap7bO2nQQNX574KPjG
w7cXkci+1LkQn0BTLycUvCFeHZT2qKfZbGXOyTBlc9JRxz8RXrcIaZHoDSkyqxx5Hr36U9ckoPGD
AFpn4Zpqz7omzpPjekpsRedWg78YRNOcSumdGe5X7f8pn94RBx0ezyURCpRtv/LvUX/KBi6LuUGS
1Bqxhv9Il5ZGJ2ys9CnieFwYtEKxbbd7RqjwSCTmBNEx2gzxgH27wizNjREXken0LMj8HEHHzIdB
PNKsejcDoR0mwN4m1mQjOdKm/Hx273v1FrHdWOdr/qX9xUl2a++p1xX4JdQ+e29CWqxcXpl7482Q
NYVxzHRthOq0rd2erWMPVCv4D1Bv3fTSRszbY8gt0Ct2DClRKdcmFklOdfsWkoDe3vbDr/C3ccjp
Y5QD+EzdhufKRgnzumG9R1h31kEuSgkBoIn8Gi//d4e0/wcjpgs4riOehFavvqchUEeoDMr7Xx1u
rhDxhFNyGxYIWY5W9MEUQZUPHlrDe/K5bHj/slfY9G7s/1j2qPN74f+4LRtHrHnFI3LQWUyrkvU8
P7PfWxIfbJFHF3ntEGXIjMMblJGIS+FJBcKHifY8IbEqr80BUjsGiHRgd3j2K5udh6aHAh8JkZqS
vZz8HinOKWzM4+tPWHdZ95vWg68PP1mFf+D7WNsBJ9s87tSmj1GP1kazId8aw+SZV+wU3Hm71OFp
ot6+DHU2inhNZHwoxefm+qYn3bBfdLf7+KBe8hA8xQJh8wtKgUG4v7JfyuvEugHe6JdHdgitXd2h
ywfUcolNgbsysJPZZBzFpCRC3BawgHtfE6P6OMjO+ZyAUNU5og9sCWAy6Vook37O0Vctt/epFwah
B43J1Ecm9tq3HjdpdQHW7k1OO/U5x3JVXFYArrxbjSY7cJwEyq/DPNsIYG5dsaujGyK9FyMM3qkw
LaW3/Itzxk926YBWI9Xy/DraYbI9Y4uj1v69D8Ddg/bVvubjX6jTZ6RnRkU6ElfEwPnXJ9+gO0XS
/bvMlAuD8kaArQLjPeRkqd5UBnWaGH/qpculZ4Hs/nIHQ5n/qeQOGPVKvJv/SBrZzpWJM77fodPA
XvHIFJUKGXTurHFWUOgAxSKCydfRYUpNT0mVllPz9cICNMsvPhV9Oc6XosGtVETyD4jKxqIGYJEJ
L2YKS+yVx5vR8ScG+03CSMvnTI5I94H77IXJlsMNhD/gpyl1h8KlEivTyOMjjeJMVb9asZUN+My5
eA2EmgkaskGaIwE8n1ICkwN/K0c9V8aT7fpOj2AwLjR0ei79b80MbHyQHUiORHFwmsAAxJ/cAXtX
vYs20H0IWQ02m4d82ICacTas6J36W2zMMhPl/vp6gDYr0ZKMwFErVzRmRenVltlvxtrdsjXR5MML
7UNFkl1gac4nDfo8a4WMB3HrLnNskncYJCMX7boP8pBQMIydX4T3p8lunAKvPwJRrFd0bAyl9P0B
CNwFbQzIvmByCSDMrnU4py/o7HujTpS7yXhBSdNI089VxKeaG0WwIIdp0oDbBDiPIPu2bPuWyAFW
9y3L1GFYOAhSHiInFV4bFn2E3N28iqOEfINNDHfVn45NoFVPehQNrLgKYDlWR3sISS1hWkFSHWbh
A3/mKPkf1BKyHAyutLJgtWctTg6yOUkAUWSjQTDKkeWwDa+yRmPjXGD6JV0vHvwNjWMGDAVBJmP1
pm0AP/8jXWkhfE1U9/ZTwz8HUrkPPd/Dy8tto/YD32HO6pmx/rcbETcbs1BjLICMRIBOcj6MC5dg
+QLl7jahEsIDIASqlQrTauJU8PkAw1KO7C6VAylGmsIEB7SuTdGH4AAB/2JxYDYGkQ7TBf8L18BX
LuM++mbrJMEQmKE9v7Kudhg1Xl4wCBEPsFnZcKaLC7tED8CdDNetbZ78oibZEliQ2UR59o1Aw6yo
BOazYMBbSPh1HBEPg8iLoILZKLRDsmvQ4DAHFD4v+N96NEAj3JezDDipvgyvVlPb2jqeja7GxvE5
DWwl4lCYmFuXj87hewQmC5r+7PY5LWCrWkP/qmc0J1pk2q+NFzr8bb74Gh4BEDQYQYFNDjxU4jsF
qewIoYgWVbFv2Yoa9fnVCabP+Z/KQ814Qd9k/Kqos1t2MeMKcPpwz5Nyl7olWFN79RxN8VB4Dpmg
HnSwSepFo2pggK3wSofl5Pu9qgmllPW/B/zoNKkuZ7sjtwYDJt5aUIoOVEBL2Eq4nTEe+TSANqsm
ZaFnj6YbiS1+Lq3cKix6mARvLpcHlqXy5Zh9OJSvNABF4XCDw28kCNqM6KrDpCpkQNvjhycL5zCx
qTuk02BLNuaM/fThVfA+kmwXgDYObsd927F3GhrvzgvASt02AGO5D1UJ8VzspicEn0D/ywZ9NDlA
xm7JMd/S7IivkgWmcUw/RGzjjPpx+X5VlYgFEYJ9mu2XW27zm1OCqigG0V4+OQW6V12YQnk3vyNs
XQk5qS6be8Sm8J9Lyijje5hXxxID4iPaIkzgep1a2tSz3PIxFdys484zr4aHYXjSIL9yn4q/gEMa
gDknFgkh75ap9naA7F9K2FEDtpHwdNrzr8oX5kxmj3K2uZWgB8qMy4W9ydXTbymozsNZthH5Q9s3
dZpeELSGUXD+VDVBIkYUu528cwJCmU669Rphi7NWX5BCiY3bEw5TfNFxBTy5ipPVz5mfZwfFJ7VZ
FXKeBC5vJ+lbeZS0xEk/qoAjJDG0N8XyOK55vTCybuZvfFW7yF1Fi6C12TAToO6Qt/jcnCRsEzJf
L8W2eYQPTYyvM+HFUR+hC7ASojGGRjfqs1ZlEMkBhfI3nFyO0RyUaUP0l2kTjPOl1uVjVPDsnt1p
JEJWt8xnOij/SSR/MrNKluFSbTh8+RiLLI7r0R4j9dUtilvCibVQvEqtOyrretzearkHef/+MXcz
7nH91JElt2h6we8zyfIiVG3gVhFhUQO6XwdsOSuhD1mjX3vTa+6GA5xcP2Q78WKq0j26L9BuhAnD
14TU8ZF4jVZz6vR8mUhfeNhtDE2ouAsgoKi4l/AQdAW3kKfN9TmeGcQ9ybznPud+mlx5YXy0lPk4
YVSzjjcIAfpFAkkaEQNPNKHG1XjYZGyFv+h1eZv/qErNayG6TUm3Q0F9frGwjNXEuV4Per0NwzHU
dOAhJoRuJWkvfUmLDorZuO4qShgJdeLxktCihIQXxTH8UELHa5n6k7mx5r02+GaKOKFFooWQ3iJV
g4zWKZQBg4roRgVi/APMyEhvb2cccE9SAqVHHkTENucAbG4qe8hWzEVwfOURBJLnJe6FnNaq+oOO
HbN5CGZxKsK74B8bmlZIVIDn4bs/g7ASnW/vc82Bn5dKh9ww5yTLsn1TTwA11NtOpGVodLlOHcw+
JCa1ensLzSfKlSAWZvKOdMkOWcLvvn9QHGocyhXhmfzrYfmXnxzOFWE7NVqRfPZbWHHfYnJ9S0VX
ORJycwTgtwISBRvwY967QkCE/pD+t0KpI3qplMuraVTe0X1WucMJpSbyIuN639MOsVGk0X+RVVRo
qSlGWzXUNHImapbXSFFVoilvbT+GFnyv+2OSL2exZZ69bz7Ec5O/Trasyh9UZbBii+Q/vs6a9/uV
ydVnu/V5U+oaTVh5pT7QdmovY5DKYUfHzxuscfT8Wafhpn2M+SUwdBFpFPSXxReRj1Wdbw3b5RPL
HTa4c0zyC9qjx35XNizO7WUV9hh9wmflYp/9oAjT1jovmZ4JPs5jxLZ5ohMlyhKd3njx0hWKwoIt
zsp3dcMcod9/PJif7vnLlR+8LDxl96eV7qT2NXaOEoHiVWd3juOVEbtJ+owMqnpSRDQtWQNaoxiS
aloUrfpUxynjLZay2L8fh/Gku8G5olxulfhGtDE+kWiJzrX08DTp9BAAY4/d+MvgfpogWBcQDAss
0St0TMGjWclIALS14nzZQhGOR/ypGVNaX4MaovZCVfeQlfb6lVNpVcErYYOeDvqbhW00GOrxj3ye
ATdYoO6fk5HFg5I+0Dty0cWVJFhsbXm+trcLEjoteVDOYpW9U6OyPNamcQiiQiEIuwRim71zyiqP
Ws/WHCsREexaNq0D9YpjlUdlta262cLSWsi5zdNqlk1m+MWNeixm5wlf+XOxlDBs3BW/VxBO4Pwk
obLoukK47cunwsodApeDd5jbZIMDUi9wZ5gr6RJACTuMzCptQ43tUM+hkpqWPzCdYamF/+h6xad8
6hm+gQ9Wn9qL+PF0ooVoHBan8nOWSknY3fNLu+FXa7S0rlW9cReNCONEOtSAI8HOC/s/LaUUjiHB
lRQwsnj6ITwNgTkgNzRTpJj7htd1TcmOAByoc9AOVUBPBk2ZJC1LwAOTiY2R3O+VfhqjhhKp5mN/
9eK+XJV0YjSQSLRyCvocBASc8XZXihmUq0KT0s8gbnQc9pfjFEzDi3ak1CUEhaJgQZaYgmKHK8rP
/5s6vpXlTYtE7iHRDFIxr0ZeYw/50gw1OhyeCrlJNt/HJzZinIcKXWrKIJSEFVS0w5kvZK3Yl7b6
xNf2Eionyxu8/z/pkhgmgezMd6wqfHwku+5d58MHCDRObJtkz0lSWtSi0BdG2k1WpWWzsXZuyu6S
X21s+i0za4xBSbeZ8gul7KpKW2D3fmWb03NgDL5HDVXw9+UvD7d9q0geAT4fQzyg7cBX/cVLXdP9
SEVNLTzk/ActwZ8vRkWwnJTyFuJ5NHGdtwWmThO7sUOSVUd7HBhDUBE9oCcf8Yixb7eNJEDYsPLV
+cwu5eo7ZMJuP7E7HR0CIT5z6b9DFDvYfBFCMugT71WDL0KDfVEgr4li6X/wEbGS3OQ0tQSh/bXC
iDJOj22X9TouPdQlQzR0Do2sV/s5TtztIeZDh5RqZWgxTObEJpkbMLjKU4Q1yvJdmfoOqGl0yhuH
NFMEyJhfsGd8gmAmWeY1ymOXZTt1qpW6bCvr0GJDkKZyJqfXJm3dkau0MA7lpFE2XXjhHAE5QqOX
s+xjYS8PvVFMQujV9WWeFrKJyw3Yc134EMu4aDSS7Ay0aW9ZgQtkLOolgevC0objFI7aVCuLijW/
x5O5eTxfoxLpqqvMO3GVteQxynjq2Bqb0YIFQqTIeMbbMAsG72q8jgIO65UvRUzFkO1/f/FzC69f
mJajjUC6EF6DdKCiBYhDRA/HCWYQWbFpEMva/PHzNZyNDrD1196dR81ETNPONWkCl5vkQWkNJpUG
y2fzBUyi+xkKfhYK+7TOWWsKumGDBkhik9+UpPtpP3uV4WIsa/2HzyH3mlnRh+kJEGPpK++0rKNd
YZ1vKF7WsqwpH/bYTRAWhvkusJgD2pDLbSxA7oI0ORWvPLOQ5ZeRL+4YYmg46SVvq2l5rWyWUVSb
0FpkMmoU/EaeiPHLiM2d96gb4D+LhspogrPuXkPYLOwqyrqzDQTgSD2b+vbya6nyYuEeWPc7PQBT
1WlxJfNXfcfYqAlAVD93erJCPgRI+SVwul3cP44LkHVBFFiNQz1KQLP8bpjxMUYITv/6RbQaMfrL
w6Ef4S7PI5/i4n9G3Bu3sEl72s/4MykoHLDkYxxpZb2Egf66cVDZf2nEXU6MZbY23xaiH5d7tnKg
vMVLJP7qSGG9L9Jg1ru3NFzQXs1o5m37iWlX2lBVdSLi7Y7kTUaJB931x+00CLrqtMbzSnD0GsTf
v+g3VXyPgIeZ0n+amxOZggSkJf/SMgZVk40OhfLjdxY+E/Vwfd7CUScvEetDU0iauL2JsbiWyWGl
IbLBbvNirSCNKcXPS6DHCAVN3KPTmxW1zhHKvw9tIVdEeBTetpJrE2quV2CTt8xR6BufF5vrcyB/
pzylDQD4LxvzsWK2rF4ZdGYIl41FG9iuxs2rofjLpcyhfuJf+aMIudPbZ9Nkdt7Qc87ay7PI7jmo
h8yL/DNbwY+unBiq/SPzqp1ydRHlHN6r57Akvd1cAL2PnNjENCk7iEiJAbCx65HTanwsuW2IjMDs
BvAPe8TSGly+yDXnpwTq6S6HQHCDV0rnlF9ajQkZOeITTLV9NjYafyJCN3fom/g4GzMJDAKNzUeZ
5zFu2KgcpZAEeJu7LMEfEZU1p0qXH83VSCm0/8Qg/R5I/obIFBDSMmDo2kMFZ5lH7U/GtqDV/7B2
pBNkgAfsFiZ7IknvKH+jEcHXu+yyNcTRhX4GQxLljQ9sRtuFsBxenblgCwQAWK6yFNRrLYCXiU1l
0qO/ie4d0jXGAxe/dNyuQrD9lWTeUJ/P8bQtno4Rc3iqQvH2+UCRP3+e2XqueZUzi9YXkxi7BD/G
gkpypZzUjBcatsW/yoHvL38QIYlfCImCYgejw9bH6tOwW7CnhN5Z4bnvQJipAyUNRxjB9M87tvmr
SXCK7pf4mnMUovEGUa5T2ojLAU2o+MFVFsCI+F++Ua3dogazxDKLRnZseZS9aYsvIUs3BQ6NDaC2
ZvWXU/nBjqLOhNB4OnsHUweVXPV/je9SgHVBrBMgSm318T2nw4w4wqvAMW+8ISwq/kXHw9qiss5X
WSDXUxyp+nbWGPF6W+BA5Xc187InZc1uoDZGkqIupDbBkKys02tzzCANenXJTUtO0isSoF1M9g8o
xwo8fJ6BiF/VCJg8LwEvuos1Wz0zciO44FZM3nk/o9vXUsk2YE01KhnN/0LMHXtR+m4QjWg2JeNc
w5ImKTCkwaemtVvO4Ff5U2qWA29hsCPv4a/3uS5xS6lCyT8WPz/4V8uJNY2gWfZkHtwVrexAEa20
pYoA5dUc/3DOghoJAlDG7NYmf/Pl3yFnj6tDyZlxlBFjazc2/pbt8RaE73AKpp97JosWQ7bovgzS
MCVwTNjoBEaRHI2YBiIMAZFAexqjnAlNMsF/wxlZNjeOG/dnqrVvJIte/A9PB8oQzO++5ldiB4Mx
vYCdjo3RQ6qrSzFPpIvy02WPDFAgLx4WxitrnbFs09RdPvxOs5MFaj6CTZ03vGbb2FPD3zRpppVk
2WBoGJXv6zuwH9lZ6ZHQ960w891aiMdsLa900yiBO8ofcYuS46V9xEKISlE0G5ThSa0uzM+c27o2
qLmsSPEWTLGbfDKFFaOxcYHn/plCjAnNnztyDwN/EFYHrtA8y9Ocmu5haP6I/tYx1cLHLMteTPGW
3frpfaDYc+ctEcNlBOdRdK5n/0035Zgi7olGGV5O778N2mwIQm7CZKzoE3odOemEGNd0szHyR2xP
GrjFqFKeap80PrjQsZw7U/1Cq2Je11r4+cA9XXAqaThbVzIPnjSEjkljeB4RKxqu/BVOv/1Ddmio
hdrnnHo7RaFkRLZvEaUJv2reZgqQynk/76lwFI2JApQv8D+siR8MCotHQefVf+SmzAkuThK5itvz
8CCDVe0hbjykP+az0u7duJ/3asezxPVbBIUtyKhmAmHsTiLg1SQL3gHtQXznyl7F39WbGqIaYdRK
RpwRhVO44LfiAqt0w7V5pRN5AdwlFriR3/IlnqT0q+2kEXCPqk7SzEjV5zpMqBYlGEJ1WMeGSviT
zZZzf1KwyG5y5EeEtAR6OTFRafgwNlWWgM88GaJy0UZ+yJXoTfa0EyAjm1UApkDG0jvv1Ttki+TM
UNHcmzEpyZjZVuo8jo0B3/tXn62LBoqTBIERWX0UoZ/qVYicD9DAOUOBFurtIKiNlCxawWxr+8p2
ksDstaU6/GNIdJX4uJbNkSiuTspfFueoEP3wvcyyXfj1OlVDFzj+mBQlIuqEdOf5ZRKhiyhVTAvj
leA1EMtt3luXgIlifxmlLrWx7faxUP+GLM18C3v8CBQEFKRoP3N8A9/bGJgBLBuBm3MgrYkRRdJF
Zc5jUZ4b+ZK1E/HdsCS1cVy3xM5yLQSCCu+UvzSHL1dXA+iggteTK1+9DR/Pm6kcM/ZkBmmkd1dJ
Dc3k6ekI9XYJH4AX1CnSVjdNFRQE3KreKzk8t8ehpGZ1cLPiOP6xvVGgYTYMkGkt9p2eUye9pzgd
fZJQEqB+HOSGEaxX9baYdVAte6IXyy0dIw8TZSH5zGkxWY5TjB/bI97v3K2cJadgIsQutKbTwKtR
HIlAaxmVg0JOfj6XkwCA5Fz9wu9ElpfDsxQRv/3dG0rmzTc8TZZyB3MQVOeOLtu0TfprUfS5cqDy
v9eJV69j5cZgt1xyrnIbDf23XHixeWHV0Px6UxlDaFRutMTcldENpzAAbzzsJq2m8D6itNRc2CuV
jOQppznp+fDRFK8CTjQhjGOS9B7qTVzchHjRsBLHEbCnvARWCN+hqbGPoqo4ZKjSJk+uqze4Prk9
6wPHLXMQJzVouELfqvdIVM76781V8CDdjMXNIZlZBMQtjPbCWkcCY8VzYI7dsS1lMoAz65tisMXG
X6VAjI4ydRLNS/Ii75WRiMeoNshNzHBZXvAPzSCnFpo/kQJz+m2JiJq9oMzE5B0yMvFRjuvIJQ+B
bH9SSnQ1p7/Bs4HJyirVNB5a3LjqPRbbHfEJv5dmqH+3HXaWWO848zye+/ju8kPZmRQpeUagpQAt
Rnp0gqSL5pJU9NzU25jn2K/VWx4CTG5BLbSh8LXszydI6YKdXaeTrDL7egVPCEphjytrsU148YUG
qDc7evqNuPC3E6QDZZXHdW9gh5aeyR5vCz19aAvqcZg5BojaoyloPpzKAfY/Oy483I1ZHETZlA72
tLumSoTO+ObLP8VkMBlaly7GXIMInUvkDoCsPjVRProq7hdzseLWDukF4069Z3JV7hU2dQo6yCg2
/lCqnWfdifmxzZhH5uw9ebtEXtUiXO9qRWGVsVKU+WOPOu2dD5DwFuXehoZ9UGGnrW56fE9rHyea
wGA3VAD/4yvySAmHWBjcOw61DiLmjD/olUo3TXRsgIToSAgOHDTjgmvcJIBPiywv/N58qrruSjr5
DSIbzW0IPGJqPscwRb/6fWpuQfAAfUVqyYsiGHBc0tyPGQgkSxfqexD7UaG9r16AIcpOZIO9vNIO
BUxgawACUgb872/3pxnJJ2zO/F0ykEpA5A/9wXzDlDzMJSCRPwtQynkSPV2YI8xM+WgEDWxygAtW
DGgQaKgbZwWfyU3BsA5/VhMVPEfkpWU5QncAZqaYCzFeW6Oc7lnAxy0IqNIOSqMEIJ/HOZRfyUWd
tpHhLTDRCt3E/3btvSicA6H2V+M/DlGshpeCCq1v68ky+Gs6OsSnKVhlo6EwR75BnL6rC2GGB/M5
xixyn2RQPqDvYg5sg8b3NnCRNyk8NzOKMtZ9d6AMtlEDIs3elozJMVLXOpZCKde05rKN6gyYzQNy
dxZ6854YSSnnbmpt0FziqAU37nDrW6uWWWfz1k90y177jpu/0EVL20UGegMmvMZMEHv7bBdLMnTv
W5vB/gUtTD85pl7t94iwNM8900q0KcYYddhhKpW2hw1K4VbKw3Bpnz6qX0/fU6amt8vbwUPJrAl0
VCxxcQNMszGH6amBiit/DN0Tf7OpfpFikt6Dr02f9NTaYAkgbUKV4REl7wLEBXXQjDsoKvwKxPIp
RfFHIFQ9qo24FSW3KHGOD+5UexBjFcYDL1rsS74GRsAcVFYPyYRP99iDykvGc3SDgeMd21l/4Z7D
MX1IwmUZOXTxvNh+Vvl8zEaMzP6dNprnmo9TclvYZRgbCVJnHG8O5caMH32mwi65TsTj1fmmbvIG
rGPAMhWdV09keDCVmB6Y39mpbaxo62VtOd1Hp13ONMqL/i3xIChQCg4PYQYMf1qLF38UC2bSmhdb
UXABT5k3my3HBQ0ItDJPPSQLFK7lY8xrHyFhAz0OHmP2YEoQkQlTPobACSvatesR3UsyywgO/Rd0
3uIr8XF5e6RTvnbDqHJP3mmPhiBtym8lcZi8Hse38pqQ26hbs+phpDQHSO6xqON0aMFH+NeXemDM
0a4geNYksPQ6aCJ2wSsGp/CDSFHdq0j+BcXgDWiHINd6mC0VtzVYbNI0sV89mnLYMRUdQT1BAzcZ
6ecvPfYGhLuV2mQnLp5nFilp7hQLjkolFz7QEfuUehWByayC9JlikLvlP5vTtK+gr5KFwWV50ki0
cRAkVOpJbya4qCcnSL1TOEQmcNSnsJoNZZBMkJyP27bf8OXw7Qu1DlZnkGsrgCfxTDYMWxlwW/WT
QbWhlcbijQzKacQ9WTepuDfNhb1g77VcTsjXIn0txpi5Qxdh1FKFWnWaZJp+nuxBO76OfVqMDd0S
p6ecRxVITjqCqSaxPnNLETANMSlwRE/+zvpOMWhpUC/0Yu2MhPFYcwzcRI7jlE0a49xKkQie3H2k
xbdRWcnOHyNajuzEZDyHuL5jaXrtPmG5Mv4GFM8TpZwDKaFE3JD7+ELWwFRSoJ5O+/Ni/EZRDHRU
u3/QjVqozTIGQTw13sI+5+2Iyc6MlWGj7D1t3GtyI543THRBXM/deHKk7aVYm0100pk/WjQY6abm
5ZVTdruvdS/MsFA1NbmWBD8/TySffqiEa+FKhFsSQtO5L24+N/uhf9MU/eMVKknuMBA/S/rP1RqB
8KRWsuMfh+1zGqObc/rV8x5A1trzOy7NrCxO3/l7b3iSdpCftMMXW09Dva4ocsDxalC2vbbRv4AJ
EBs3Db077KhNhFiwn+oqYek07lgY8qKVUDekqPTDOxwzwS0CJvblV3AYKXwaY/lmkqc5yxD6eaIH
/OXUAV4UkysaKtN1bbe17h7iVCXipHc8MVahxA+kOvpRJOxopWuqTxKUh80i8cweZuzbDN1J5tBP
o97NaS9qS0pOvG2hb3WINjbshfH4IfN7tL69/kdfEyOOKioDKvYus3CyXzUvlNjcT/R6Ow2wREOt
7aFM9xw8ItGbdlPPVKDF+8VYp63ikZhbLgrqmPSM9HsZCJLAzHuxm/HOIS6K+VKn+xwD0Hpdgm5e
lSBUNM2eIjYGNru4rtbD6LtpDNKpLFtXlhQkxnhkM8s3bvDIq+SjQoKIqcH17XPw7VyNNBfd7jrq
o/sVezhObDuiwaTqGPPEQyaozBX4wF70uSG7TC8mCAXQJN0ZZ9PX2CkTeT8YmrIp6bWAxyCuhudR
SQUBp1AJiz+YUGVvhiq2hKQLr76vwNLtmj3jCceYOr9V1vVBfZk3d1suesz24MgSHFKJFcAz4BdG
owp9tbROkGkudaX5jqFVJYXfsiSttEA7AvEA9e5ncY9TNYSMVYFjYwmdhQEDZnCDP5h07NXIB0g7
c6H66r/RPS8+rVOe4KyU1xJ96z5YwzRFfJLAV7tE1Uy4/VkUCumPXJ6tm2Kye+RMekcY2vIMYRCY
4dJ2MsQlGGOKXBPxMk0RpyagyMuaLRKfqRDJV/k8OTNmoe0Nv3/CG68z4S7bxj28NHhbFSh1C+y+
ux7YYWS89j63GxztCRnjCdxjtyYJMTo+LkqRh6BvNdR4qNXgL75OhVvfuo/DlYMEsByg7MT1PvM/
ffdecuJ2/WhaoPUeiLzKtQKx9fKSOs//PcVWwNvtCeWQ0xV2mKhK4nK+O+mKpe0N89VI6/Onwrka
ZnlaYAHVfSyzKV0CWdN3b6NiwjFZfeQhejFr502naCaqYlzk2CLOOjhXYjBUt3vpe3soazjwrrv0
n5qP2rYPgpVjWQbyuTt+urJ+VZjM51rEZj6dpuYLmEC2epUrEqrMKGfFemxdyD/Jdk3Uv7AfExzQ
T+gEOECD7JRig46MGCA8i9OU7BeNm9pVpgqvZ/f/AzX+GX8JeBGnJBycmozTYzxpmJazOOYi6Si7
1GLRHmK/JMuAC3+ILtFgA4BjeFhA4mHFkqArPtc7/qscmZwIZx6+YTMjDF2bmuFNqne8zRula/M4
8e3FJfF6tfZ6GGUKJrs/Zh941LqUnj2wWnstNbamdnYcInB30AkPaR/KQJDWHENjB1pYGeXokYAH
7PS225onGjdXIiV3tZmUO0OHctkz6gjCet7wiWLnmclBNk96jf2UXs/dIvipEbgtiu8pDo+D9ayf
VfJRDfxcey18npQ9/p46i5XJqLfJyZod3RJHz/kKKxtIUGD+u5vpLvI/YY3qvRprLHDVol/GrhAj
l0z6gj7Xc2PUhOQDIbnqftkA3VZe2mhlO99GS1a7kW9MisT7ZkeqF6tsJbmcuOid7vOEZUSpeTHu
UIZpOhntmTVVV7S0SWLzNsJEgcjLA2uaVUy43S8tuqGzJTMmTmgAByBrNX2ex5FXdsN91zq0mp6T
S8BMDmajIZmc5ja0Njuy85+k6hVLqmtiZk4r45S3f3LZ87wN0ASFR5VhF4TUjJNirzwkceAwUoW2
oKObRrDSfX8ASw7MkwMbbQbOD0ND0xxd4WaUfCsfBt5NAnigoD7sm4qkLdLYY3336vG7LPJTGFgl
CwjyibrNjojPZC1w0/hNgPqS2hf8OndkpDoYJO0Onv/zsXNwWjvTqD0eqjqVZMkXTXPDBRT+ON1y
iKHGVlIENdNkQGi10ZavcNZ3OSvIsJFVrEKZHzFvZO3zQR5N4dqI27eoqPjGMN17IT2ddkzrO39J
pTCgEU/RrG2YeX7nfj0PfWbJRpJvB9TxpHkoLY8gWQUL0z1ce25i1FMKc0+pJi6BnsCPm7By/gMn
2jpRljbfLomR7abUhWSBZeRKeFwYRhce1PZwqe60ukf4XA4Ndg5216Qybg4Yq6JgJTUbtRFEYWQz
1qtpg9jXtcartPY/CiMKfRXLKMOWDTDAaqvkXicj0AAinDwyKV7tj1KvGG9rZRDyy+dvNKkCmMDj
eDptAWxe2zCZZUuepfxPnBVKnCmAMi7GxIYE5J5ryxZtp6mPRZiVKo1mQVn9eNn3vX9+4uVqd/VP
xa/aCPZZWHM4tPju6Gsc8Nxq7AgeM2KoxuzNEmVJ9VARU7AfKDnFFPhDq6KTz0FMF7pn090YZ4Lz
YItZP30XPfG1ycKT+GOaq6ERNkFQOk2z550N0T/tOFopXzknymTt2aK306dD4t91ScIqi99Ulll6
uDzbWqbuDg72dY5YnGoEJnGMXYr+9ctxPgKcZfUSGsEaqiitLLSX8QSChltPMdTywHEh8+eXPIyR
pK25PQHjMfVYEdvfL2EPfre/L+hRlxyD/KKBBrY3DtuvKbT0O0yhI69M1Hre1N0xCzlw3aV9DAst
WEMXLzA91YOezcFo2VRPG6uVwgkqoNnb2MB7ZIbgRRuTPcXgFyRv3jOa4f3CTygRROrXrtyTcxM4
CNUMcBsF6I5JcLPa+4YN+wdOe7D0nNK+NTNyyGWbFz0NLzQIJ5zetnq8pdtDe5MqeJqoHT/kyUN1
IsyXa2ARoSfjZGprhrnZTJbAU5PSj2Si/IcmvyXidixxaiTjTR2Yj8SqjR29WiHk1KPaMFEjHolL
3vaL+w39fVxg+xPAJs9gXlBdha6THJ8NdJmDcCIQHYrK38dxbbYLcsMj8ygfVCfz2/IxZ8oGvrSq
Byaz8E9vMg8PvYNJZA+844pQRpREtTYiXtSmAKOpcqU72Cg3Bpy4NlGdlNHPspHwaY53H9MeXIbo
/REojM+TpDQCa4yUw0KPlgw3xAfK0KLiHXG2C6cKjV5kXJmt+7M9cjA0JXp9zdIsWp4Hc6DPuYBf
dp7GSmyNJlbFUejJ+6AGgIAEEh0CTEewpH1Rn+l+JqqcszLeLrKp6SEZqIIeqVneuVMO3PtRaoev
mIRJPWpBQtObJDuWt06GGkz4ngeRQUjllNNyv3RYEi21cOSzE7C5FkQ+LVUHaYYHV1oRvvJLqh/E
8b7brn822RypKxwDCXhJtUa1xNnLL1HHc0/aJbhPsLv2cns6uJUziFpz/dtbaUDIQszSDJ0S66lT
BhgQiLgKEFtqReoIFXg9mHgHBGL8i9DYvuE7Td+quokJwh6amSnFHLtE//7e/VTko9FCAP07T8CK
H/f8uUpJTYy4vOnNIp5qDGJ1BeCt/Om5Ni4uSZ26h3it4hvrcVhE1m0xXjwoI0bpXdHeH0C4D1tA
BU7/YAcuOz/ocbrw1O2Yw2HQVEBZYtnP66QrCiyWQtIQCXQ96iU3/R9YgvL8vUDu5AjI+my+GD0n
K9ztMq2v/PHMo7MUzrJWi98djXz27iMDjQlwjDK8Tx7o2ruWDzotVaPEojkbpAuFpFP6LmNFmJ1S
IW+Sb2PT+UwoE7gP6TsmkpsNecx3bfxbJIvUS842uucnhEBjoIhtEXynePtYvPluNg5Qc1tyGPgX
qgHeIJGRDMkrdPeu2k21+b+FZazZPPYNldTY4p8UQVF3kR3lmqPDviafuZh+UqWBqhFJNDDvgf5t
nmt8wAubNQ5MXf+97S79nEl+hHn3CWNdQNIk79sR6nmLQINX6CzNB1+9tkQ9K+8o/fcrPvi2e32J
2qdZhAerGlZAFy6q9xBLGx3oY1+nKd2KQ5+N5xQIiKMfAuod9afJOAZR0olqlkhfW/aVaTAwpkZy
+6+RQpmzUBPDGn2l8+wP4+xbIVK5U4NYtIbYVdAlq3qZ4xYErreuBBC3Ykkhqt3BNIFX6IbXLlrG
MMQcDVVGoWNuriKGNJZLIbL5VPhEmzvl8NWv3mRMVNmgCXCmigW9cS4Q/Rt9iyht73OjBKUFJ0CC
H+NqkaIVjpcLNGto1vNRqOBOzn1jjxT86WXNBobSxiKuPVm/S+Os5Y24dNwAo9dC8VrUKlvsmQp9
trfQaj8/wMaRB8GOvP+6pists3/lfeegY9uBfh79XCOM6zDw4BUQWCEWumidm4c1a56Zflm46ghi
pdpYD6Rrj82tcz6nC9yoNt0NBYXgMcYQJ8lO1QeI8r9XXsG/bnAtQ5i6NTHH89C2UI6dCrEqaD+7
e462M7jOLJManw5Vkq3jFfqwD/EIdo3EHi8LfVBpBEGwEbAGhrVML61dwQayP0hyrrChhjpKJJIp
JRKICZDxqo7//gXvsTrDsKUjqQMzsZ01brUQcTbVno1RkC9Ih1VShT0ICcAFlt7qbQO+CPEEz4kW
wjuIbto+lwGKrmcpKe9Z45p2q+4/5+YyX7ArcvhP3xKd+Uu8xtJeh0dUhDHsQtnQVbsgOVvorBiF
Tir8R9NP3rhqRqpi/TujX64R7tpsfDTARihfIYqErqm57+KArYA1y7S6ZjB/gVkVTZ16w79BOXLy
cMwJKcmUCGczcwgMbD7FrZiX39lKfE0RcPxV0WKkSIK5d9o65hzJT3AOsvwrb1Ft+DZeSkolOOBH
C6d6U1kP7sXpppiRC5AS6URIhEAooOxffqtrjHmrOXvpuIJLWetIZNiNRF3TpDBbR/ZbrmfEXBeF
JWp9IaVyu5tfpGtsKZf3tqG/rc1bH05T5173wtZfNjGdYgsQ24xGmJKpBJISXTuPJdwNYo3zRVSf
c+Mb8JQziBDOuNnowjfiAFk5SBZAo9IltqmxS6gCF1h9aJBGJTSrhPzoOZmnoSjdogp2MDCZEbVI
gqFBBHD5fEygEru+4NBH6BKE/F0VzjczK9JUb1wbndQ4fadN8dBBGRmUYra6FZF4A+xMyqHfCgY7
Vve4RGyFP+ecsJxpHJACY+m8QE75pHRYSVDp2P3QaZQrRLewdRqhxzULlL6ARinKnFV0aV9tNWyl
8amUmwcQScTOsDsBU0KQfjSbpKukoF7ZsfRt05D5PXiHqEZy6JZ/2WnIPIA/s8GSCC0qxKICoU7S
5xAQD+D4hgwgnDUW+zAzn7Jk8txq59oulMgVh7a5eEMWzOVnebXCmdu2J2Z/09N0SywuMFHpsfN0
Eg+6tOxoyFSHTnb3K2up1PzvGlvY6KMIHnyuHaZBO4tBQCKYyWYPG+tDTc8+jKbLvyh0p4sExGn1
CsLRFNlpD35uHuHIVVRaYHB+Q4TVkHArtM3QXCtoTM3YpgfukXKfJ8FWyjHrNSGXz+che50cpLPP
hb6soqqhV0QqUY/LDJiDX0nN6pcdusVs2+nMMUuB7PlHc122wrNR20dkOnXwGV1u2qcgrd43tyMg
OJF4/nXHIVv2TkARd3xBBdQpncXvCyJMIUmhQmzsi+F9xOqMlxLW4Lmju/xiwBisM9KA137Qni05
B8d41NWmB+9OX1ipAHVdiYUW8J8vt8YdmHe9nyA2tjWE5fPgeJc6SXuPG5FEgmw1+8JAMY0KcVkQ
dC0DDHYUNClU/n0zOZFGT8A86EPllgVy8sY3WkNqVqre8hF/fDQIXC7fzN64i152Cg5mEPnuD9SK
/aqJT2SU3sJjfHH4EwpkuW6baWy1qMVrToZyuLHVNvLXp/EbD9abyiGjBUdkpOQQ4wSZyPrW/0jH
xVZF1OLVoLBrI4pQmNonQKQZ3xsEGOI9SEjm/Yy3Cmujvjx6NZxbSWGjBd+RqF04tvkBuBxFGuZM
BqSbERjDnh02qkkf/lkstPkVydIqO5a10rAWZ1/hmll3maybChWYa6QuCMSHSP8QTxN2oV4Z/KGD
lputLoKD5MoqKlNqRfaXjA/Hz+O8uHCxtKN/BKsJIup7aUiGlWbNj4GUjcOXqt+4i4lJIUuuXG6g
pMpPmVmjoakrCUHadmIFCiiDkb+2+gOtLCwdM85JNB8kdCpdpMS6sQ+RqpTDkhSUTnDrKbcKT1kF
+/hWMEGbGy9+RjHE9WxRwaOnBA8dFr87Dce/qkDWLbet4Y+t5gNNy7rsMnaMfNyq2oTWaaqiqv5z
ZfJ88OFwE9pXJVdj4jcvOwt46aJROSdgvkO4h2uDNQ7zfGjKF8gGf33MJPi/e/xsW+3bav0FmxDb
BR3ycp4X20JpWFkoO2awF8Zwlxgbsad0Z6Jn4FEW1uHk8V1xLlst2LyU39TpVrS9uGV6QNTsbTtI
9LzGlrLNmgr0cUuN3uFry18yEdZR8Tj7l4Q5NOzT+iiPfWAoAMs/41dIN/I4vXkLAAm4zI6R5wDS
D+chQ+6VynmF1C8IpXHr43sNgE3x4Wj0JH01EL1pU+TCMr2PkrclakcNJ2rwLlUk0srSqe7xsXZR
Y7RvjezD46fz/1y/RAi6e88BoGqItaZi+wd7HfDgCYbOMMRsBf/ywNARosOQx8GNhrVT1TkmGxoh
PhEx8f9R44FxvIYfbpTx7vMtbnSZCtLyFpIH0MYbGYMwzs8TOyFVFptiW5emzQcWeR6nFuRmtHnf
QEqtiyxd2sePymIl5T8q51trtgsdV8aHDcUIv3gDaoZvOMqH2d2YWAXIMsJZnylFLJApSsw0CBIH
PVDug9FmfIN0bHt8iQJMQYeJ23H2aUR6YppVaCfSfDODj7WOEFQ7k6khloQOW9u9JiIGYFqGaiAm
P8gqgeuLmbgEJgGIS04072B/On5YPEyj8EtvLJ3Ufz2bM6l49OtWiZL3ua3I9IiMUZZbJgqh3Uw2
57LfWj4xjAqk5ceXRIbLVPX1OlYA4g5m/5b9kW+bH1Eo0Zpnd65C2fCl42Qac7vUshKAc58PRYoj
BRVYVERTtHoJlUIpgmUmKbIayzD6MYu3lReSEwfiv9G0YqTRJDL+CIKpCUGowWrRU+wnEvu7hz7C
lRZ8dDRfQZXg/l6IQpOvu/MFVO3bbVxmB5VZ1g5Ca4Ucj+ODbLJLr+8kusy2/X4HZNyLts/sfEmN
DEY66stN6rR1XQVhc11Sr0Ez5D0Wr1tidzwgdKMNnudDXZUJPQMFoirfQONbWHia7kLQvLIIjiij
X4cKZGiKvQgRHrdd4Lc0WIIWgEcGXUDeWEVQjlVdX6Ff2n6IBRFgFxfxDVoamw/XvtUVZD8EIsxW
SkEKp7ZJAzoGhTNEO9KubUZs8F8aRqGg+aa0iBHTZ31M/cL31czPYXGlGjg17kI9k0IpBQzclNqX
BLzH1nIf7Wv9jignSQyvkALa3y84Mx8noxMT4Ob4X8thfxI8y6Wh0yuWpTeaoKgoaf5v+9f0XKqz
v5IUW53xxO4QORaoX9IePQIrOnxYY2DWCzsibWJmGGhVPl6wHHwmvqXQ1+UaSMyKd+NI/GREwDlN
7qMzpDrfejL0L8OGo7yClaJp28SbY+pjov1+gAiQMMkAFGz+Gr9diQ9yfGzZwchGOcYGexg/lsLq
j8Mv7iCOVrfFN069g/iwpq2Fy7du/Ery1Z6bXmoBodQDj/X69drC0sm+EbDikEVzz0adpZxlL4AU
7VP0KZO9ptP53r8p4lqgOptJKfNayoO57M1qAslh1kwQZ9l1YmXp2GHzmUwBV0rVrMreMPe226C5
JDxIRXOwz9jahwuaJLyN0Cwm5sVguqe2294NSPmAch/6eFbcXUQ3TDwXTrirRdq6PDL7kamIlJFx
H88ikIvYjuFetBvpPims75fuHrcxlPMkEBnwO+kk8walT5QVWuPWA1P/3OoNEmGW55RfBxRR21W3
qyKA6JU/Ppp6rS84FHwV+ZENN+EXMToysyKfLO8iiuifHvDcRvwra2HvkfkhpDA70vJ1sG6b98QG
raICz2hfnSC5JAC78Ng2uPfBJ8G42pNyWuHItRElZ5JoVnnBgQg8SwbSXZA1Hj64+ucow759o9nV
rjVyvVYBp+RIBt7F3XWbAEvOzRZCeeT/aMyOSWHMKGXTfK4GGZwNMQJJn21gAg1ME89I77aFZHRe
gFaJxX7+qf+y0c4nYPdyQmB6VKA6Vdc+LtliJqVFWQoZuW76nLMUB9BgM+pGAo/3YmipOktd8MT+
t2BTBgyV1dBI/S+jnDexsCIFcKmhAXQM4AIv+syNgdkXDGJCj71c/aK6fmJ1BX9Mr51aM0pd1QQ0
i+1hHUyRVgl9wsvhpxhjmS6rIAit6ET8eWlJh/30QCZVKs/LIbz5/n3Nm98ZlNCgzIWQhhOjY6EP
9oDfuYZvamyDniNjSKJix8fft6Hf75AozVRSJ0/a9cm/U0P0ShcqrlDREA5yceMeRQpTQ93/RZU4
kJYk9SZj3zTM3BT/QDF41bEdp8AVFyP9qB0joOOpUg9WRjyXPA25e/edafSkVzqppRtB0YEz3pQF
7VlM6eV0ltWs19ZYzH6VXjx1HtsvgVZAOhbLUQx96f8+W/dmbWgt9bljkrXBM9TqZYSxWmgyloHh
1XcC6+ayN0wGCE/l8Jzn9ozpBLRpDDm/F2YWU9xL+/QmenSeYfKQct5S05Yaj944RC40QnNOtrum
52zqYsFIhcfEZjhYrZ2j6WAk/ZpA+nLSIabDiKmLWw9K8VMz8mPxxje6RAR/tEfJqk4jwPSR85vH
xbIn1ED83UqTw8uw40ERo155gcMIbBELvLb6oFtZYW5am0xEVzaT+5BPehEV7jcaBuI7aHIx+fEu
dC29zrZVY56G6vE7HdSdhIZgZDBYi+36TRfZpkA3VPbulRtd1DlxGKklbqeiIh/h9jiFPDOp3Wuj
Em4kquLX8WV4XtUBPaOKUfQAXoFrIzDWuHU0ND/MoZtH8A3wcV7sPFCtCDtGSZuCqJLpSGQgXtbK
WnWm+7XS++9sACYMgEtzhSiPPnADX2FqQ8cdscMDB0VUhBdtd2WFIqM/SobU5s7SCuNpwIKKy4Kc
5CqnkuZHi0+Kl5UBc3PnjAuIw+riZJyLuZuzmaBr3lAqF5fj7XhO+dNizlzd8iOXEtSVFem30/6N
kPwVPjx0uBRp+kptCj1hi1saWqAcF2IeqPKVd4p9io1siL2/TyfBBEdSghZU3xSGC19nauaCdubD
YbUm+NrYWKGmM+nf5T+XN4rnFbFxSzWOQvoLaWiOv9H7EQ6UvPmJOq0FK5jXXF36LgJE77LtZa9s
7AooWhXQOYrGRIjmzbGGqdKFKPCiadj8SjxrqERmwI8pg+S0/d6Oppgpv5HQe+xbHocJnZQZ17nh
Obos9IziCcSf08cmS0Krhewx9deSEuSJ88I8gjru+6btDh4nDXSdA9re9Q5ZPnetOCiEAwmBY59H
uQHTQcU4ssLVd21w6N6akTYpUat/eN6n64TRYv/Nu5uq/OjFVG/EZ/ibY2VQ3ihNHRQUmnkI7i4h
Y78+okgcQon5dwdS1ZZk9bccoja/glSExfIMW5c4NTia9w64OW6OsF3kI7EmrUFq6AG4chnIq6wG
bhMP1lRZoNRhtrHAoSF09uAns6X/C5TCBLJx2NsTO8YkxxoXsbMjjtdAt3cRM8WIlr2IoXPcP+yD
/FzpuMjD6cCVLcX1zyTUEkHeTe8J7dgNhq9DGO1M1JVB0LaJcQ8AFVJIGWnUvZEnusJUW1o6Qt7x
cbCv6lw/gZPJpQ28nmt0rRiY9cMbYZMIcLQ1UpWtKXlch5LrdCjXN3z7DF8eSzdHBtKzJBjGwiYu
j9aBP6N2iFTSSyzNIoZ5aM0wvEfVSEWHZQmGWfgra2qvekoH3sp5Az0NbEFSzKRzZO2UE4Ap4oNd
VfmrOxW75SQuCGurlc3fJCsODLDIXviNRKkzZ3Ifi4sW03J6NGbXLbHyRif6oC20N8UkTIaybggN
BfemdGqSKVQ8dhzIFqNWfY/sSGuRDh0QU5g9rAGtALiqY5Bact1iXxUzXgW/e/Or9Ce/oYwiIlwS
oSqUZFDQYKa5beW7UIH+VRQwHEpentBrLtiJk4TL7XknCAVdi4bzrLHOwukkxq1u/qIziICnKMpR
WRWHnD1xZDp1De44IslwHAJqxQKFsYnp0FKsCzHyOQrTu6v7OgGSGcjb0y2jHqeRBcLdcVSgXh7a
iGmklkI3OTNYX0vqDoWOfP9nVSi7SfS/i8oTCULmw/3q3KyygPIeQvfIsmaLClMju5xOhFbDxQ+1
QvF9USsPB8wMDlOP1AouyXAnUitb3hQ2zgff4ABQijZo08I8IZI0VT/UKwMKJ0Qf/n3XnYELWZxl
lnP2YRTN48HQwdEy+gJGTjTNZ9B8d5/bQVXyg4LMP5njdkH4HF+4URwer+3qBidltEhiFT08WLAw
FJK9jqReCPxiXNpUqw3XZCHBCuCqGfFCgHNKLQiPw5Tz1NSS1ozfmKT3+cilforKTv6RBsvv9jRb
drVjh3XqMWv60EV84eMv1FH3PIRGq5/ztzgDkFZzT5GZtj1+IMQKYvem2906/jcIaKyaOWzkj1+a
0c0o32smq+Y3oaCq/+MnDNdb0uWlXnNB7BLuvOcqUTXdQzC5OvqhidN0cxAZ+yyx1V6eAJHCLnFv
1K8oLSWF8l1cntXYW52BLkLDOw9efhCsukyf5ZMV+IrxHt4MKHHun8krftChQlYfV4Oc7SlmC3Mb
Mif+HrKNXyM/uUDZ29Yye8lWMhbbA4eo4bokQRWEuL529XGRhbCP+1IdE/wACGOFdi99iBtvFRrB
BCrgNIOUrL5Rw3jpEx+RAq7F0Ld94FtsrmzMpmZTMZWDhh1jaW8k5MnxXjCQ+0XCOMkU3AKSDFi3
DQztPrO75u0Fz43UTFiuNuz5oaKuo2I2nnImKlFCoUrA/B62X6boXM7GZME+bKyFLbpT2shgX5Af
edp5n92EWb49Z2K2YJMqmqkxhiFM4HfP44Rpz9QbjKT3xi+uJqRoB964+SPZ3fCjifIP04oG5kf8
yXxAT6O6gHpgSiFLah25q2+nCOCaeHbuq4oyx7WrUf+7/80IJJUrif8ok9tYqFVuaV2ICqqdWE0/
qD7p4LebTM4tRJKUj2DPYcZqXYhfM+TGDGa/HQ9cqvNhHk7KbHhUrfvXY8xEGYg3yycctikDYVog
Kq8IRXouCY+AF9QL4E/3xMorHNQgUO6FmNaeAsQTRkfn16LjKrEVmoVyALkXxE7em40czZ9yfKai
VZYGDIAod/QaEerNPY+a70K8s5estzwDiMAiN+utfTc+2nCqqriCAPBA7eyIgGKV1SY54ONe4lBJ
PGTiaRsJzy+DKkloKrDCz3eFe1dtP6L1EBkqWIjNsPiz9GYHSrqH7zRYcG1udL8Fhb7Rh5d3QtP/
FdkOcoR7prHwZAYH0KnoBHf4oCqA+fNgV7CfehQhdJht0nEHB1U5xpR3iKr1i6YTRpcL2GPs4NLF
btPtUxAWVu2ePuUldRnKNHAAqgD8ICKRIYPUv12X5vu5e34UP3JrYwbHzMdZ0XirVugkG015u9Bx
G+xCynL5K7YHSPI4YzsSjsS/LiNAcv4TbNh4UWy8SKpy504f9CudbPbVBZOXDypqBEgNYMSaE3lP
pohGlPPT4/6sQSrm+NRmE4oZRDC2wzbddWDeP8nqSj2hP0Y7Ofk6J72JJRep86fd4NrJCla+fXr7
JfN0LGfv9r0kfVMD+7vGVxyWqlWwK+KzawCoIJEZ1B9FlfAfRVSkqUn0abNeQPA18tUdVuK+ZVEv
m6ceLYCjf5UgTKECKjsP68wxVuNfXCB8p+huU/ZY2I1zOxobP3vBA33Mb7+qpQUOze4QFXkMnYBB
AImcrJG6FvAUBhjPUhQFEuZQodj4bXNUgn2wAWvTHlxvdgV+DX7b8I8vAC8TZlY3Zl4AhpSrt8uV
KnJrmcwCUuKs66f9EofQH8fIlw7mGT1f+oFwkw/Qwsnv6XaUb7c/kRkMY4A+JqtypnvBtuUJUPgg
8tePTsC15fp9nNTzImVArCmcAOVU2E7BLkj69ZJA0zEUHVc1DQirimxm8YfDpoFfFW50QxRzaM/t
1+Mdx2zw3BVs4bFhdFSFGG/IDTTxUXLWQ4hSlxBfHlZwEluJjlwjnBeymnNgY8Hf3D5eTiqdAQRE
ggSU3xWz3YouONnXHZGYYg6InjfCeR1nwifh3Gc7ROktMn7kTw93XPfXhY9mhr9gnMe1ztXKXjfE
rkrqwYyyZPQrCM7HiuGCkMjL63nfp821RrErT+4CLNmkT+WR6T622bVWrTIE7xmT/0uvdo5XU4Ks
MOIGxnjKxvNqcvKqWiTHdUTOAFa786S2z4+6nmb+ao1LOTbMlZSAmIASEsI0ieEoWEPI9KQR+Wuv
fQs+fR3bdn1qG8SlpbudLa3sHRfZL8YS50SR7liG0Sq/PYDIeW1OpVU9Fs2SFQh4US9leWWoyLip
C2VUjWKdaP47Iahnxx+ytjq0MsSP9MeUPPiWVwI0dMDeFCs8iMh+aIM+u37BIugIbfDu0bt/6s8P
O/jLTK5rbHc2TnSfnC7XWNODwM240BKhB09XjYFgUmscPc7m+lvtFyPqk4e0Yc2k17CpWqGmx+8u
SehTCFxtGshRlh67a6WVQp9qKBQypelezi4OR0krYMEN7zgDu8Un9fvlxipFOHo6y477ZtzNcrUN
Nrlfm/ozJ2QSxla9QFNE0GA0fHVEbDmrrM4GoVoBjDzKdw4BejvaSdzerSFa8zAYCWHtOGC8Vg/P
C5tq3A8QaFAvj2sR5PdCqmMnek7uFyaacG8Srmn0eRNAWMhEO869tZ0bODYuM4SAgwKrlPk8y/ve
a/Qi6QUeRE+9N1v2BhqZKxstukXT1QUrSg2m4NjqOt3Gww8oFNKurI5ClmA5rJdglKVCy3xGsfqz
LjVPUxdZrw6d93YRpuyYmNTsDXOf4t5Zhjkm16B1kOMhTtRKLqBTQnIoCOwbcMlvx+aZkuN4Gbom
/WV3kWVrVg8rDyonaW7wN8GFtjwxb/P3NWTjen/hHW8yH8IYebHGyUrSfnOs2P3PAZRzIx24CTQ5
TQUgVfFbIg34x4sB6DdH453vYL3KdBcWn8aSbTSo8BDpGc3WbqkjATScS/8VlOsXFSegwQNU83Yi
8kr7V2oOuV04Qa0ipd2AQXFYMjaW8pZDwxMbRicx2d9+8sHK1tyupdHfwipp5HrkD5sVm8aNonJW
zlfs0w/Ee3Em5LaowxHtH0iPZXaLN4W34Vi5AQ4yHnfBHE3lK+M7aQpkpJJG8OfjysXaYEbfKhH+
eg8ReT1Ka/kI0KtR6gky5ztOOv/Fw1cm0T/hDAJjEQ/mtwMI3m/985urGtoaqGGdqQ99XYxOhuiJ
WiS9ka4bxkRjJaN9PndGIla4IdErpa8ori1nLz7xP5PKdnetLr2kPodYht7nDCm2qbALoRAhJqlp
7aUcLxPPmeUjpXuiV/CS7MOMsGUbqFD1Js7JIqUQaBpQc2yjbacfgxn0BaazliuLMlEv4MTQdBAB
SBrWF+OhBpei5a+2IiVJhm7hCwxKlXH47vw0MbaQjiYbcSMSAUGZ4fG1G/Ui0EjSB3EpssdcspLW
6Kla1NoxdxmOtqjWzi0NrJxK+2NmyXCcQwkAtbKs6H0lMEkfN9gKZKNRu9IDVMxiRXFXAUWAEJTp
dfFrJDfprqUkTPvUwNExOf9jM5D6cky658kRXuluE04YWLbGoUTfcj/sg4PBJ7Z9ogBkCjbepJwS
P+G5DVWjrIRXHAHPwdDqvHvqbLqIqCT17Vaktb4Cy66tr+fAPK4MbnFgflabsfa+nO+CV99DRpXL
06BbeAfRUUKrNy/Q+B0ssARxFRNYoDU4xG5DWYjdK0aQv8cEXl7cGCmWhf/KWioL5ke6tJ2JnX24
O3wQtfH5auYty2R808tM9VvA+fdoSX3Hw0/KcEo/yWxObYWC79kiouFsj7qG2nShHIuZK4SAeQB+
ybJ9/02yohGJXYm7AlQzmEn3TPgDmYS83G2Gj1SM7CGj+05bp43mPoOMCXvNDiRKXdQ83SZLHqoX
oFNkjkCS30lbwFcHiCSdxEk4irS2sn+nzF/Rr3dz98+fdJ/lebhQRiS0DmEOjf/KoTZb8dLA4h0Q
MYG58SeR8mjJM2DjrdiP2QdpN9WyqmAVIfN8fatJ2WiLQMvSldu9La2Q7SGmc7ruDnZMf5UNVWw4
OeYtEEDgOyGdqvXQpa4IKBnYuexWZhfxwopFoMYjn6s5EHVKRj9u7KLEGEHMWDnlqTfv1Oq/qq6B
nFsGrz6H5bS8qw1IUoHwu03vsl5bvaZJSgxHsGhKCJVaq79zQtNS2JOa+9CVrJ/AJ9qdygx288LH
yU42RUpI0lLUByA9ES1PhreVXPvJRN6t4lLTQBfDu5T7Wwg99ay8+Trpc9bdPKC8IZDFETLx/a0I
F0yGYxtXA+7vCUGkavyzopiUbEAuQ7kxk5P2miCtC8jxRSZ7yHIkHHnBmftenjl1KOtTq75NMSB6
rh9WOywI0ZFgdFGAwdeKgRH/n5zkgWmQFo+6LZ6SNydsb+WF6bIxjQRqxnavjQU7YI49jfz85HtU
BV0cQ+c3zYnf8XNu4HhZwk7TTtdN0Ap5cNEyNGuSm2f/VCnUiUCglfn8JvbrXsOIJnjkgo+fy6Wy
CJPmxIkqbzJi653om1OMZIATwdNweyHmGbo1V9ujX8ARVDJmt/3DQiuPhLppSonFjiANf3tME/Oi
B3K1G6N6Lg+xv82TTfMKnTqufCsoTMhVn7feZ/T3VLQy51y5Fkk6KAE7gyNMzUffDf/+nYt9yeX3
nvooSSIrdCv7NB5+JyLT7cK7PfC3CgPU9GLYATrFKVEJsWTHsYqVjh4C5YWyzJkp+HDHicT0jN66
rcRozp5BkxWXdSKkTqZMvFtfgrk4oRcRMW2zVZmw81r+RZ1XGVuJoBRwu51wBRHlUVF/NyaBQT2/
6p/Fxu9iGljFtKocyjzlfw/DZU7G5RXEkKYTwm2I8LcIzgJTVwNraTtuBB2YfRV3hCpgGUcR3roe
i+R+Si0IfgQL2aEEMvTJxr62IdiqY0EuBqesD+5NzEifNCZD/iEWHmVxk6AThqK0YFqGG/WKWAXe
Qnb0iAl3+sZoIU0b24jYDZX+d25Eb8lLG8LWLeVfP6H2M6exM0gBNzu4tR7E1pQez/8fyGJzb6f3
cF9CxuMt1Ane9VKQFvq9Yp5o/oyi6q05ShEHfex27cKvhnDHQzZfJcrFRPSopOtpOCLW21P740jO
u/gajl2okRElcg65Bgd//hZa5WT/6c74immwkJunpl7V7CDJr20DAthF3XFei4HuobVPXUx78TSD
AHx9qF35ERyvZ1KMPvhS+oXMzbH1N3I/67lKjsh3WzhUOrWNzR7vASLqQ7U69qIHX/sOSH4EY6hs
35I/v+2YuBzhy9oi38HahvHR/2DctzIMrxoOAZN+k76Qsbl+EDI7eIwLBJROhHz2F8IZ23SjP7Z4
sqsawqrd4rLJW/JeC6AFquEeNTH9yc4sELqJPpqCwa5+2Sr+qElSlPp5gZKrDkkmJrswR09Dbvpa
JrLnbN/igD5pIiCo3g7ck/nSfMoL7b2EJG31N3kiSTG52PjMjjtyV0o2TCnHkCzsZmMEGNANkLDW
RlOT2hQzNKJ77FRtyOYKUchM8fO/XpeynV2tPcy1n7DSh1MUbRq/2ZYkIIOmNZWe2cYyFBfrAReP
2vUM2HMOFYXBjxo4UvcnL75nF9Han2+vgeMp2WiCVrOn8lYpESUG4a4eDchUBNg5DL0ISd0Qnhwt
Y5kSpBsQ9qruJbbe5O8COSBaPD4ZmUpPKoQ8kg9KV4dLkFPmSpNFzHt/JiMHteijkYmbxALQmg5R
B/FvW8V98ylqxl2udQlMKc8q7oH+e+Obi5khVZ4U9QhKjTB7IusCgssrwW7CSUc5QPB00H0tlQxd
uqolv4PNsvovOctxVlzxJyjDlNELe9YsG/s2Q3fgOFyRIaHjo9yUfgamQTGNIEFmq78z68eiGFf4
X92HfyzHMa9vV+uItvFH9mu+pALfzBpYwOsOUT22mNoISI5LGq4uhBPUNrQAPJqPHsINOBHG0m1m
ykVYzhrczB1MhE2pyg8W1epL0/IPhbbH/+9nAenZLxtBtibmp2t6Pjzrv1t+6U4hTuEjeoa3UtLc
BYiR6X7XOROglGH+4DGeIYg3NIjuf7BPFuOEbE6CaJW5e1H9UPqDAk4U2kzljkvDiTYdQ599aQKF
TBRH6sOiIz0Gkiv6SY1PqGndieM1ZygnZ2+NZMBTdZI9bKTDyXVOLTYeqvCmWYgCZZ6VkJm5u7fR
nPpNMGl6GaXtseAsflkJUZ/97k6lFo7+w3+zUkrmiBydjHRgTcS/voQ1tcvctWzpNd5ocY5bwf7+
QVKaQ404p2ACZ3HT4I7Rz2S8yfyc2IFVkSAjUsI0xHEhiYmdUKtKA+Tj+0ybxJkjLl6QfcJvm4Jc
6LCMLM60mZwdbqYtebVbWjIx3rCO8OADIrU36QmtnzyjW4DIKt+RxsCtFUC1noe+LO7P8hPRhqvl
iss+7oZesqI+OesO5nLhFsmUtYgAAGsA3EmViWmle7Qs8iF1BbAThQKkmQkMvfv93iU7qKZo3q7g
MYEw7DzLQqGWQNxzVWKEPcgzkb6tLVmwZcOrv/Tz9c/eM0CCXTKqGaYxNstQaCC1YYSGmxpU7/jf
IDpBmTsO6cR/Dv0ujzFAqjS4pMkdhP7NwAwM3pEzDCijawZyXllouL3YzwcuYf6rPUjKm8WRM3SX
IZIa2Qy62yVGxMjm/G1qnLFL+0ntYLnG8cO1hcIQOieecziX9LUF7Dxc9ZDjoKv2hUQe+AJiGdtS
liTsHr3Wlshj03xemO5f7dFFeywTL5lHRS49LUtDvOBNCsY1sDB03nZ0iPgY3KWrNnapC2368GcH
aNYqp/kOoVW/4p/xnJwjYVV+81hSyfbJOz2BC+CDu8s6+K+2UeamXuMMC27ezhA2c1CDMmfk3jHA
oTuwFchBs/bulf8gJO4f8HAWpzl/ZmFWcYtBX1/BzjnBBHgaSKUKQ/SR5vvBygch4fcNcIw0Kxjm
CC56/TGxLN68plmSnbdsLQALubmbeUBAgDn1/jveJEhc/W2GAtuUmmzXe1ViYBg10Gqnlbbay1Z1
FFiE2p+s/X4NO9dCIUr3vy51pN+t3Vabv4WwNtL5yPURIuVOfu7CxuB42YD/a8hSxzD9YUkdgMrH
lmzLmsBuoPohyQ+ugMsNXzMw+vF14n5Rqlutzi2NCr+NnaKVzjS8EMg28tYWmecVAxzGYQWhrFIG
Qv2yn4F+mXYT0pqKxtgwklSLG2Q/jjHIqMX/+//871hZb2rlruTugOZMuiWlHnZVBn3j9mxlyHXX
wV0ZSB8feq/caIH1XWJn3SlLcg5AN5KSyVnu2pPAYcIvkFlJ0Yg+CzY4PUK9HoytFIpkuAgqRJnc
jPZw92Hc+315dDRtSipJsbVmD35yq3Z/C2zTaA01c8/AXoWBYbWfl/aObAxrSzm3erhG1D12H9/P
t8zHjYcn6Y0MAdvy6FY46hRc39miZ+kiaoBAhp7fTrNmFP+Sq8U0wjM2UyLwKralrLEnggcgKqzh
/WvqhhU2Wfb/OlJqnyPXoqQjdKJdUly5m6ST+zPSJdTwKOU26ApArqxeDfR0bSFXOJdEITNxMOoz
Zz5h4oOH10n4hGoXy8svQ4997enLk8JWi/w85G2G75fI31FFNJfno7nEQ739oWhGBASk60iUhSlY
6VIkZtnGoc4EtQOIgIgc9I6vRUnR2jF/IM25sWRD3zfbBCxfm1OCa8ux6DHE13hmzftfyNvQIkgI
mtGfpU1/s4+X8eH23D+dYQS7ONFBLwwRStLpPhuXGuLcoWhQ0UiIrb3ATMuUTuKinHnwnGqDzjco
WOVAiVzuqDKnO8LzvnS0J+B3IVMxXr+TKPjhpKGVKrAE7/yG0ZuKFgTtPBaNVHisIvsmvM2GXmpa
hNDueSzLnXqUJtGU8Iu9mJ1JC9jGGbjFt3bZ7pUpBfCdwqr/mot6T4awXE7mLjpRq3Akajk//fd1
6qLgDXvbynRnrq/FzHcR9PDqCzw5O2/RAUTSJ67xjz5L+eCI2V88bvruIxTdUnwEizyxWqjdkHLN
gzJIf2JEQcPCmEKV7x8gtr+PG4UPqK6AJ59ssVsrEFfH6Pk6/bk+ZwxJC84MFcQYatPwHZyFbpsn
ratLMQXlpNFqHSGXMscUaUKFmv+4/CSs3V1E2ebWeoEMt8mXa3Z73BMDhOzgZuHW2srmDasp985x
s/rLVL5lBIpEUzGaCraXwaWsezfQJJJnJFD8uScOKLgcPpmbQECqxQfVytW+1AVv4HqmV4j84uKZ
B80aQlX2Ld9kJ2A5PIAmtOpJqLM1v00d2Yni5g1Hj6SGXwTTt2ltMwZeTwz/c4lQcyiIDFgKGKNZ
t/fJv7n62Cq7t6hywnJLSwBGHml+ACgsUHLll0AmLAgUSyIku8PRP9XhrZw+GkhXOFh9yufrxQ5U
Z1OmBAdLBVDIHbSSCQjw3pgVYmajzVQZH5P41n0ScCqEEw+xazeZwpkNAhjVvSdRAdg7CBfkRmsm
qOeqi+Uh1/0rGRms6KCsw2CmPoX65nzNc5AgjEvnViyzoCJzbDio5GPFkGSv0ygxWsjpbrFRboio
ZgMiwHOtUvox0DdqZQS4ZfpwoejH7QN82eGHmmBmQtbpMaIXt6aSxhT1MUuS90wDi7//RanTdCS0
CjEysH+iamheZjBTUBQQqNZiCXMkzTxqURp7KwUfT0SvgWi+loL+hIIpLe+gnp6aKRXl7sn17k1x
/menFxP1sUTkpW74rFZ4LEvz1+BiUtGbGKEVC8HlEu7hIUMVQzhPOlEtXPv73pSBK6THZlDGSK7d
fXw4MvfvvLoZdZl1vNzEuhZdAwzanVcTGFwGuFrjg13UhizIRCnQzV6b01dABoR58TU9CXzmJWxR
DW/44QHFbQD6z1YBWRJs3medxbTbQL9hTCAqAwmxW2+a1HJhOY+Et/NGTxAbTgehzKQUIIcx4nor
iopBz8cviviWGhAGsdkr65k+5NeKl8FwlWyJmpYUobK/EEQQXCiKr57CWc8S+QYJJtoLfbrdRDnp
wZR444RbB+yhCAEnXqi71CP+Z/TLgplIhAN2BBwhK1BJkl9m9wzF9Kkhw1/YPblJ3Wg4FSgxaLIy
GLStFaGNrpiR6HWp/APTnuR3JHvoUe4vUdNN4g2cv0vf0AlOVOlpwjoqZx4pnbxj6hDAW2v8ksgL
QQSWcIvSpfaRbFyF+kVM1fEf7sQ59LqPO76C1cR95mqBAVt4EL0RI6psVPaKhMjT0ICwzRGDRyH7
1+iOwU8+4GRFZo/YtJpFh3SfpHVoB0wYlWQ9wyh4kDm/+TCuLRB9jCGxT4zTv38LouxV0smuIKLX
hW2oSdC0Ydn4Eojqz0eraDSdyQPyFpws9WFNAl7s1N0pKP4E0bK4vybz5uYzPpj+SyCwrwDsZAQa
0lU+gmcfCfR5YggztXmRJ9T2C3nro+Or3dvTMNanp0hNUgRdEc3Xda7e29X2M2DluADwn/GlSDqQ
vkzlMYk7zquH3nEWClqeJPH6gaAwVdhdP4E8lm5XZrkFEV0D+VyDfpBShKwEeX6NtsXe5N7JmaSI
Tpwp5K3n1MKppQLpRfavikXjF6thK+Hr2AZIZupDX7AHB/RRqaqvZyjBmNulrFjzVsdm1EnuK4JF
Yc7m8Zki0RhVYM23PrZXRlJUXXZmejD9OUcaYS7g5h2cHzarlWVmJEBvwLfJ2fGEJbFQyrl7OMUv
gOZs4lCAt4I4NzfF9FAzN0lLLbmFwAJtqLSTCekMkBi462aq+1/bbeFpfSp+6duNv/JfH5kL2oIt
j9156J/RT6lMBIG3bQZcrWiiVJTevuoATTp/cDzOp7eUxsC1PIepl5NYPsO+1vZtesZbxudOcbyS
Wn7Adr3y8lPwa5TQ0MvJDBF6aumkhevVSzvK80Rz6lYsNnRhnfSZyG66oY+YLR3MxCZoYoK03xhZ
DEbbkFSKuURwyKoGc3Fkaxq9pkP5jzAoPr5Clwk2tZyuKumonN2jvTdvBtNsmOeHlx/pQ6JhLYPn
IiddtdGYf61TcfVj06xJV+byAfYrB8uAGZlJTj7RXKj6l+1NwUYca49UomiSojmp4xmJDhLlW03J
Hgjut3tcXeKKHy5BSIjdHhzx31W2NFgXn+md/6odjYk7S/6Db2qyYFspqFoB8gDt9Y6NNfSm3Mc8
yuO4/8v6M53y7f1aAFZ2tI2/qKlCs32yTByPbJAeUH28+jAfKc82FVgbxxzJGCBf0pf8EXR+tmgm
Qr+PFP5q3U4dhZbqodQVSp1uYkkjAg3zBrrv58w1GXd4JY6mhNbG4iJ3Yk6Xo87vDrou6r+QpDKV
l2YqyIcygMzDgwAlePfpGetmPLFQwL6BmT//rfcnOCbnEgnh9JR/Rg1rbsCT1WxgztCQkpW4O3c6
kA7/1KCJL6L9gsxXZ8R2oI6LJPjgxVzOitOxNQB23kt6EfAoZTdREGoKSB63Ru6n1YQxBTtpComp
BiIi7ud2HSns42d4ABLM5Uu3y3DjinHPjsKPr88V3+RsBpnKJk8CtjviXbkDhx0bHkx3CStrqFkK
JmQ42TnFZjp8hFjUrpahysSPpoF8zggIxFhD5mLUJGhCm3MtQUaIuTqiEk23NNi1fuiHWnCfYHId
xsXFdlJtl+0RBFCT3qFUEF8YTOIDFvfVdNfnqNx0jmotn6PqdtG3p3aiP1rbKpn4MyAzg6rCh+C2
c9Cvkire1d/xqNeYGu4m+UilDTGMyoqIL6VcL67nk+HEw82E9MjB9poGgCScC6zCr2GJ7cC80Syy
g2iqN4IOCRD9b2wAN3kx+1bPzbiI9C4BZ2yM1kupTMpY6GgFR4CcrBJHZu5CdA9ozHgSE5BdRN5t
Q83mzxaBA19xQ5Ci8fTQsXV/JD61MCrIwCyK/Oss101EOt+80wuP/WXZ3IJOAsu2R2Apxh7as369
x/XdXv48afZz7gSeWA+Q7XaELUjf8Iqz1OFKUAOaiYOMSNjU7XA97bYjeS6DV/KJXFYqTvh+Ppu2
gqqELHIBcVA/G1hjzyIqATLZa3El77MZNhMJDNu00Sd+0uaQpnrl/sYFSmgBuwRD0HVzYRFtY9uf
F+ThsVx8eivGgol/T7ySp85AV9L5T5xZ3qeY/wnfSXZjvJIzfOwOzfAODVC67JI2roiMW82j16/Y
ynjFmxyIfQGdp5JKg/k5XafzKOpl/I9+GNgNuIY0n/08nHkaEQTmLme7pGN9SYjlUbk185olOv2g
xGl6e12+5zPlb8SuD9kzVq64kr1R+Q1JuD3I5eZi9nLq9nctmw+ktDFCx8oHoLm26B3xEqVfcnwS
GPYgWXbCZbgFvmYm1tHq8L8AoKSLJx/McBN6wjiGy+uAccJ32aiQh9J4ikOiY2d01K0CbDY0xLaA
vGywWL5qkQc78wjEaxKd5jpFhUbmTWVgpa5/2LDAIh9W6sjdiXnbBGGMcICsYkHytnBCkvTpCG4A
2bSKWtl6FpMpk5GidXlqfWETDTbhc5AW3zIGaMbnvjmEAFMIJPFRyRSYPI9wcB2AxjciWTUnyi8J
FzMqb/j9SHAWR4u9uRGJ+gYRMz91Go0LNEkXPKqE0G19tdb1xQtcDLj1+p7TdAOoDZTmvdmUBuz3
t81tEv0QUku1XMGRYs8ZCHzW9f16MkYsSdBVoxW8drE5mlN/SCeRc0OFM/3bTeW/3DqsPmh2lgvB
eLQNr3BR8t0i1wr9QjlLh9jwSJ+DTQZGn8qGPeHEc17hKoKuEDvcynGcEiZH/Y322Yo2ouVWpcaR
TOUhXVjDXaiDdaBSJll2qeUbt6xNdi70baMhk6DX5OTHjF7scQaU/WwM3qjTCYs+luI95DyKnrrS
dPO5Y1PNV9hDaMknhTAG9sjIH1jeSbKCmdjeJhIY+q2K8fFQEti4283i8sSDYv7cIg8KYFY4x/UW
kQ8MDg10kfB51ACJB0/XjhjxkspvsBmr+lmBEfeCCO8ufYmL7FVQgn4E742PS3cQVWdyAdGiYjHC
JQYbsfENJHrnXyKN2cwtQSHY7zPjd0f5Y05ufqQnyNOTs1qgtfQ1I/2V+FPfwIvrO2sSjqy68RwQ
eg+5VNse7h0Wwp+Pcmiqs2LlrMVKC0xTYT1fk+ckyVDCNWlKde19hkB14bX95+ir9duI5K3PpL3X
yNOkZl8duQTAevVMN6Rsydlp2+3eDCj9R2XwukkDoDItchkzJHRZ2x9uvfayqYVO+MWqzNw7ZzEl
yFQrM6MO8PU+2vfUj+qdwHaLsKIvD21CCkDFO2kmNSOf1ZIYZcurZLrMQBSSvbEtwAfkwt8+yxz0
kQQqb4Z45FeCB0fZiRY7dvEdKmUTivlT8Xx5BySHIDSRMTHl7l3R66hPz1I4y+jjqJkyMKoe1unp
+XKEHu483A0IwGftAaHuXzNW+6kuiivHzGkUV8FC0TAZiIzdkrY6fJN3lLQfDCBsF3T+/yYf53oc
uCSp7pTWbTn9o22aAO//BihLvWmhiagMc1FG+zSrG5KHH1LG7wy9DgZbZBDwr2h2Vc+EF6L+Bjka
S6mvcAl1Z3/WraUp02Wlb9ETDV+OQq2C34vYafsbqt90yBI181+bNyNVU0qL9swuP4fkuSFgJQj6
yRzPn2pN0tzk0SgG6/5FgOuzUEsns20B2hDntiblf98ut4RijFgZTFHzpYoucrxn04v8geop9Xk3
JHLHXKKyISqlTSQOG77TIKFgExpfdB4dNKUBP+uzhYUiFNm1FEtqdEZOdHcnemuMaordagIHGkhm
yOh1dtqLoYurB0DJYssNRukrlXWzbeZ/RzoguaDkSrCaADa5WQVBXWchq2enNZkxTdlKsJQMAqGd
xEf/FCnG19aVlRtGBD/hK7QKGFwNh3vFc74D2Egte8KrdDMqBvQaULKKC9kdCBXYa4qAuT0ZaAAu
5ewSjsGJOaAW5ciAQhsnPnB9RqY3KFGG8E31gIw3HlRwQiXzGoWFEx9uZxtW8u/WxC4RpvMf1SMC
eUjd1h5aDnzEql7o3OQzCR5iRc5YVjPYp7g99blsmo/nC/lU+YSh2YxU9USzvXbzQM7+IEw4VeZm
zCeWLyKUvh4/igPtLh0jO8wnHb9IBNOUXuVJIRRkrt3nT67eHpo4hWN1w5VbojsDeTFpCH4lLoke
ltWt069MaqQB60DBTN6avF1T7w9e2nY1mgOLd1k1QaAJkLyAjLHfZYRB9GkCntM5FQYODayJC+C5
yayCM/0ef+Bvf6PlDB2fLSBZU8fs0EG+5czntU1697tP2xqBIG7vRlunomeOS8yC2G8JXrDWdbB2
s+YgUPRI/ZyY6/i0f3IKoYg7hTBAnVXij0vmosmi2BOhW0s2jVNJDxKDXRcaQF2PIxeTfu2v38x4
Dt+BdbvxxCJzhZ4mTbQlsArbrmfnmE5iRIKJ5FszTfadS2g9/B+Om+RHST9GG33+e+9XHD4K7sDH
iM0XXXbtS9IFe2lKmSLaAalsqDKPAOkDziOySdH+ACqRkikrIvFiEkb0T0odRaMvJ7G5uKdpN9Bi
a+uQ9BaTUm1sG2mOe0wC/JQVO6llgEK0iFSnzs1mLEY9YjWaPJWZZtWU0jmIRk+YDVlGvEHJgACW
2z+8HkV0IaeX89l1c0t+nHCUYurEYzNFB+C0sKKIHWjDFKBec8un/ibaIrUquBuxvGr04PbHTP6K
3cnbbiEaoCBFABGirjX1/i1+Ncqfb890v/BBkT0a2WQTUaGJ37noiLy4rebJggwT7PXbEHU4RbmG
StvueL6E4xXv9o9Ek/uRqNC8S/01D5mctfALZHyOFAsGxJeloz1BcJKNJ+o2ki/iaGTEfA1YBxgL
0aD3KVvnfCTVxRce+BOVmHEwWgWh+DIJDZLHebLkauX06/xuNBdBru/XtWY101ErE3ivzRbHjGhu
VhaZvGjmx6rCU3wPHL8ZxGTk0mOrwDvllpt1rbJrekbEpWeBLuBrfjRP3etEddyLwvRhIDoyStTL
udx59Td+6ke9I69S1wsS4G0Ht+ZaDa7g9A24Zxige9DU9oESS+SUkGEM/k7FG/or69L0VBlysK4k
O9yzb01spOzUiiEp1mYRna0cuXN0gnmE39Rs+JkhcX8RQ67eOP2MXIv6EhMLepmQblDQxAb8M25e
a0t98uqVdYKuzYEmpFNulSwHDMImpuNeWbsIJZxUaRcd01XvJwGE6DX810Gv3fTMDLcsxsguVzF2
IA7rc3emaRC2ClmZyXdUng6lKMGJehw1/ovG094xWsiXtJpcjo+FWbPptDbp1amajTlaDx3yFjiu
J0g2KLLd8PoIXzHGP8ZFDD+LV6T5vT8AkA6oJKsjPMybN9w/eBnuc3tY+zRq7faJaAo2fWs35jWa
7MsVKmb/zF3vHkmvWZH57+9SWiC9vSTzxybwD0E/LTBkP39A3qqO1oLMR8CJgiXOtf3FjY36yjib
Hdsak1wsowpl+hah/1xVTzrosv7UbBvNcqsR0p7viSEP93hKH/KNUPJzWKXHJ+inKf8SJb3Iach8
f1IC9KXsZpGj13hW8i4BMYsdod0dLH66j+RbuaNi0pSph4OgYns9ocQYoz93JXJPtBEMDwmKcgYi
kl9HyFXUmYISsyQwQ+/Vcd10cGjPxK3e4593eOp2c2OJcN4ViK/cemL+1atrPPQ8i/6TWFPikNcy
F+DrJqKJ/imJPTOnvh8ReRe8UXBFGORFPh2pyTtyvsT8An/sbx/St+gU+BmQnEF/BOOltVE6VJCE
gH+AlUVy7ooLq8GjxrJ6t9AJa3DH7S3a3dxFnxZBI7rj2gb+NO8lFtoW5PUTf57wLY7RSQtj5GlF
7MAvfXkDrH9VnS3VnKNYbR3js9UAr+guGRkqCJYAkqOzGyLU2YeeSOPTAXyNBnodLTa2ECxV/w1u
6mXv6SEBksLzjqlTCUrhfPUdqFha8y/01wmNGTRofEArGyWssSHx9SePcOXZknnFm0NrmsuIKdW1
tyfxEULIKENhCp0Ukhf48wwJc/4C26+s2F/OnlfeshPuvf2djxXrv04s68HIG6z43xiRoqEteHli
egbc+lmrUFkgyfxD82zXlouX5hcrbd2hk6+0qV4Djfj1DhciepzZ9BF0srp8uB0PgKVh1oDlMSbj
+LGHEKjjqfp7Kgwigm1tio7P8fSaHQjQR6iY8ItmToMRx5LhEyYsdOudjRXL8RSVRGR5VYLCNLBs
TrAwBvQphRjiTCELjuYv/wtH2jPuxc2QSwA1+q0rUX+QsWvLP/jDMhONXP8ZNTmGihyU1loAZCWU
VXZ4jx51HimDCP5WCwAyLYUJ348giJ5OYcIulhbi5AN/e9RoLVIPVrD1SiEUusW+xXXwkGKMsTlc
M70T0TpNi0X0Mg2jS1lEEDspiCMwu+7/46xsKSff1hvdBegwpscpNAcabPWJqDq9jnZJq5kVdq9N
NQPgdh6aFGzfEKlBfl+FksplO2cWxdi4vHAtGpuruj1DmO1mLS/iyTSIZHFZnFJe6N9CP2sur49R
2jJoFUJSOIawmhAuPpulEb5kyN7gSmnU/ILupJbQVErzkZs9HIHVygK8cSNIV5zC40EBxeInFBuo
eGPTaqUfksEKrfnHTckoNViqLH4ADHdeR//VOLU0zAvHGbgg6/9N16+K82iDrB4QpiQXrK+O6HRE
eZMJGub612jH2SQBkOh1ImHTecgsDDg/pQz9ZoX953GEHrKb+vLlRGmKVVMHTHAmT04NdY0xgOdo
YwdAunVbKLpHh2w4dKWdrqphZN76tsBmhNrkHX8ZWnLQsF1xdHAUdB2e0JSb7l+Xl3O67d4gzHzi
tD8CjZWm3pjcvEpVXNChscJh65JJ3fyhGn/ibmHfjyiyoB1mpS4nFN3UfKUckihmvqBK8Fk2eCQ3
uM+qmpqWln6oRfGBY5NpvSL5cgzsOkyAT+Zkdit6RcEc22Cj8qc+9NWv5XPUVaXdX6BvMjl+G6uG
FkfISnNADz47z11l0nPVA5FoY8kF82ChoMjAkIUUVhShMfHY9j9c+N6n7kcaUoCUE/AYrLYPBW/p
MOkM7l5znuh6NxYqkyK8NzxFZxvBhliJEojCcXPji85E7lIZLtcEJqWt7d497pkmdVO8Dm6gk2Xk
vvp0J3CHGaPSWGONG8YLBBACoDAGyVskN61rXf2S6xug8jvNOwwaJGsvZeLfAWNMUDgt8PuNMPoD
fJhUKdNr8PJmZJQxrScswspIYeWLcPigEy/Rm9z2Su8IOlNY65XZazXrdUSIPP0gj1HHPozgPkWA
kzIR8bzeFxHkMZp8R94mFuEWwUEdif/nN+Fdm5BEDIX+6V03uAv9fkdIYaVeDE2qrevbg+KGqPUN
e4kSCIKBaeA+MRn+FbHrTHgyQjIeUs6nFAgaRltgeJLxgDC+0BkiFzdi7GrZpkD/DO9PtvxNiAp3
b8fOdziYPcWeOuHf30z/XK8eF9j8pvpL2r2Z00ByJ2c/O75ulL3irEvZSxegNvuD2YxXU+l3VpH7
6CZjXRD4vUzD5MKg2V2HoWBbNeE0PFw9Lepz+yNj6ujqhr2k7i5ft65SL0QAoEKuUN8c52sfgXDG
vtmS39xN56jt10dB3cu6pZJ32ZvAViZ61Zwkvcu0Ixmj61vAXgXTAn1vs/7eAGylYdjca3dyKVUX
pXYvnxVtzoiwncT+y4dVVQL+25kukv3B5SlDmgsBeS9a2nHXGhL560Ei+tJn8pPr02OUe5Y0/CnC
g2nzZxAmx/BS43vpGeT4fVZoJI4JOa+K2pyBwOZVpwggoCH+JIttEYyVvydEWYRAVKpVIpQrAAiY
zRLGyrNdjskzUzckH6pKCR7sFB4Bxe6y/ZlzkaqBW09EdLs+RMiJh1q8OIGi/PHJ8bRsGHa5nLaY
UJakWHLItxpTPibjVQdKoRXAr/NKIBUg5PIOye7I8i9bF9XI6JyIAHlAf3saRz5Dz6FI7qE8F+do
Y+cxhN2NNgFjhkxw8PjRG3GdC/5EwQ7x9Tqc1pG94UJ5ijjY3gzUc3p6MdH8BQed2f5rGPkXlOCC
4zwbzmLNSCWn2wj6VoyQCmpKiEGAfOPZPXt6xeCZ8TGghTXDe59Vhlp/ML1Ln7+48SIBdYBDkijf
Iata48NATo3gQKn1RCj3f1NLjXNB7BW8nOFxCwiZAYFGBrPkRJCwCFR9Z+Qa5NXvYL+q9GoiXZ6c
Y5lWM9XABbCJRv+3oL0j2ybdNQfnNSfM5N0007FCVVWpkeGufkojloA5sst+fnLQQQYQ1V6XKxwL
e16FQ47d6hNn1/c+lP2+UuFhL9A0J7OQn6FWdADflqKNpTJTOw0ZP6IcUttbnHa+GBjpZskykP1j
twQyR+8orwlVDwbzuLeSIaVIlseCJQ3aQ38AcFgZl52bjRUPBLwab30lqdPWYvuN62G/FMM03A/v
sYK8CnKIYEL7/FUaWDOtZkjhUGOenLuIYfOfrvDJw6dOesau9tRuK5xySbee7COz1zypxDY7qTQR
SybCTnmnhE28KqgH2LcYLn6kLgzoRRVvj/Wv1AQ/UW1swWGaq9SXavaagHmQC6+zxD6h/fSyStYG
kO2/0aBdXrRghHDSp4VPwGOTbQn/GsZAlL36duYEq+hVoCUY2Qa9hQ2JjbzPFkpx8v0HnSm2awrl
Pp0ZChFtSeNHxRcLG12cD0tWjETZc6w94VyU3UvajTe5eSRhqAoRbg20HuLizkbocW54TVaJwqPZ
0+Zqr5RoC2FKhcOa6QZGsTwLfEm4mDzWHwcer30/jdlDjHDFQ8w/thNydFJ1d95k6MXKK3DNTTkl
8r3xB39arv+bgHyjuXZzCmAB13VEHrKdRm+WODFF+14k4EO99eKbnbR6JwqyIvahQyVMhr01KkT7
D7SW271HHhj997s0Voq83+WrWP+QzEVZXvGXsKMAz3i6J8G44zNWVeOqW4q05z6kWU/gEjJsVcF1
vKihcY0TrOZa3BC3+f7PYCWvu94h0HGjbY3Sol9X8WD5O/zfcI3DGVZYoNpMbeeMviA5S8r9S6NS
v01Z/ZZWVoKX9XAqpVcZlUmRTopPBINwb1Y92+ZLDR4IUP0ytmR2V9UqSwH6QJjkLkmF16/LkubK
R7hspfwErsKEMb8Xvi/3BgnNlSaacdNdQM3xxoK25Q2OZ8t9mvz6i6CmENgDUe4aGvCS8cSmUiOm
/AtHpHrrk3hfuGclWr/uMelOG3gXNotqKSZvBN4vS9y0wD2cwxuNogPSlaW+waFwuHI2wvQvjps3
pWXQKeF865FcN6LhifgRlsNmQG0lUrzem3tBXjaB3qKY1p+Wf0E7MasxeB24BE9JZjuu9ihvhlqe
0S0pd1n2jdGYLn16SWbKTEMwwJh4q8fzRSY9lOyBi+lBuBfce1bd4UfvXZMK/7riYyQNJNbYrFQC
mSNPwuOQg0lNOXyjtifJJS2bDrvJjvEEpbOajT2JFmAU5yWhl29/hTwsFsJBX/fNCcXV+OR2j5Pp
MP2xxkpMrWvNAJ3J62Ooxokc17e4OMx+CaVBlJPgpsnr7QibvIJepgqsUQUBiCrTeZWw9SYfOkUI
ZVfpvtlSuLnPDYj2Vun5kQniD0Eu8PXdQElGMrDHiDQbH8IQAqVuBCEdip+5LksVtsfQ1wpud0Tx
0lM6/OJx6krqac7lm2I7giHJTlVbOlHQEO8RjhI4zXzrNf2WmWlWzlhHSIzNPuDnHkJtjCqbV0i7
WByYKAg/hZx7I/IT/vbTVqoEoAZAe9YsUNOyv2xs2SkFkV1CBDdLrSBG4rk4Jd5Jxr7BzHO86KgW
nBMC1yCdEc8fRZGLhxMbBnWquh+0y9+UR8JIek5jQAQKgke/OaSUAcHKItzd5OZYe/ldYpOfKx0w
04N4Z+YsQXXsTJE5T9rzQHP7R/JBcth2yJYc0XsTx1hhH3RidU4xwLDixmfBbvLHdUdlOEZ4gDwH
Vlei7sJdUB0sF426jO2LZUY1oWbykdQAZYB2qMM5aeRFxB+dBzzE3LMu6fzxuTFQH5zams9pVKQb
4OzMnn+cr/XZsS/xRkj0yTcFU9qSDU4jv6Rv5Wf6ULmdx4z1fOmRwQz7y6dzw8hcpnKTEHrdKZQo
Z9NqoXs7o0f+83yxZ8RVTlCpdnVDLG1QooyeZtUkiwsa5imnajzkdhgqZQJx/KypyKUosKoy8Y39
/t9AfjYisalp6kXj8gDXTO/ADUFzdWMrr8UKM6sX4lvWr+yCkcyqCfDqvjFmWYGejm7HHhNk+MVf
oagDwGdYleCXaln7GfXZHQ0dd7HjpipfksmOG5slmS4deek7GpGI20hYa0sj87VPA3ZWAAreccrX
dNCgZud9YyXaUqeVYCN+6q6rwsARMpZcnvdR6NS6Wzl5P0HN1K2rnN1mWdeM9tDvHVBXNmk69aB1
eCH7FqVp2g8KKSTC0ySa5ypal5YfK4nI9Jb2DcF/7VppF4vuSTFPIA5QkwCBMFBIurBkmujVKO2E
0Qz6hmO6tTK3HG/JgaY2RUECHywZXnKWjsK7GF7Hy8RTcclZazjwI8owUSUOERd7yQ4G++kejFBl
Jzdqn0CLfw5a5TiZ0odeEGUXuwzJ6ZDYG/Rsz+XXFKMyUaaFTBmCDdGkzeUxrmVKnzKao9shX/ai
C/RA3Kdrg2ATcxYoLZ5vdCcomnsHq/oVWjgewqmCuQtXSMqUpaFXqD7hiBHO9KzNX4XrtSv4CEBX
fMfk014tfX/0LpCwoj85ObbUzYaD35bqESW63EycnuNJ3/X271xMn+vgUxBW4Y25yxAEw+5eMVYD
tveLWHYVWzedc2JHmnDyjLm6STMA1Sf6rll0+Xrams5AuDZXM7eIhE4GnKfeskwY/ZN15wgbDGbK
MnIKkVGdrhDDaTyC9MA0dr8/r7OpMRiw0wU5YLR2vqi2m1AXodCsHlJXRKGAVUSqoluSBHBHs7AJ
96m/R8Xia4ECczZ8Rq1eEwslCrSLT+E0JIoBJ3NNRV2CsHUhJU3TSiwiUO5kdqUeP1aIewD7niGY
lBWn1YRRlQr5UKgMPxMrWuGqghQVX8ny2xZRQdT57CQEo/XZ9hR5BMsFUgn5qvIQntb33ueQdn9p
PHb17k8uI9aojVZ+f9cAYbhwS5p4YQV3dT++h5QsnFrBAjWldQoL4Ulbx+Z8OlOgK4gnCrOKUPjT
qEDEa/41ug5uHGUP8zpSeoggXz1spq53N27sobkgQVIo1QEHCflEtcZ+hBG9EYr6kjZ4PQW4K+oA
pf4Y/XYDzBPhCv48tiHYOx4Fvl9GOHpjbHBpEOWBV1sEuM6L1XOatSkcrKXQkfwxuZ5AqM/KKF6q
1P75ybkiA8bM5hdkrjoOo4itmHg3R53Y5MIiOwAurK2kPucI/Cx4GrFkqlPffocsmkfwKcapQkmu
ou9ZvF9B9dZnwUXSQIVWu6n9mBMNz49JpsQOrt2eYCVB9XZ9zENsvO2+mrL+m1LBrGRTHgj91IqL
azn1dMqWrcKBwpwb7+2EX3ex+muOqk3rYgDEybo4Qe7yPS2rkeEW1F7tkdKX5k60Vik2woghSXDS
HWL2nQrO45IkG7nY/C16EzGm7gkbWrVpOpHfSyPi2uLOrOVtnZ2u+FBla9GVsIX2D92dvOMsNtuJ
A85HJLKWusyG7dOYI5s040pMBQ17fE0+CPsIMeqOfRM7dmB2NlF+AWcU+QVtLhtgw/kml3Oc9F1m
FpdCc0a41qKrmWonU9ZobAI7p6NZk/VJ0sB5ROXyfARMJKFeTmG/vDAPUlNhS0nSXX1L14UMtqKX
vndJ20vtTZD9LeIrPG4XyuUXpKUP2aVmOhIPPZfogYrnXZfZ8mMyIl5k2YKJMRWC9Sm/GAqjEpTx
y/3TnI19j+B97/C32Q4unYA8U0q0Zp4mJEjcQpXfM/MkfW8Jh0KtEqJp7HTBssX+B1DkGP90BZYj
lUXMze6D4TQyfJv5wNJR/HTM+thqr/JKbLLY5abH/ommRcXYxRwfn5zQzuF/87P4c+gB8YzReUVm
RlWCxUELGD4hUrfg+KFFdpK8a0ZEAopEJtT5QA/aTbflV5rDpDAp/0oyAXpRmAwtPWKxyWVzCxA/
s95VkSkkWg9pK9g4w2uZoTd1BSJ0dJJt617tosDx1IyZOrTw/g1meMafgGtyXMWLnO3KpU11cxR3
BjRo5I5birQhQ6LaGVQIJOBWW7dmnl32Wa7qeChqLtjkjbwCIz1btAhti0M/PCMeLZL+Lrv4IQ8C
aw1NrlqhUtznSRQ8imusHGBMa0ovsa/jcsFtEaTt5ogvI4HY1HwLv49b7Z07XB5RacPDGw6+mvdA
H63sczKO+GlBRoYgUJxMbOHL4Gr36Dwvi7awuuvIN+TJJzzAuE8wvfguwECLUuxcL6x3ADgi5Msv
viPQ7lr47ZTZ9gi2G8F8LpCjEi7f10CzkkvXyEQ5RJDe3LXnwpARtSxvMF+koBqwjXUWYe1WgZMK
IgC4qf1JE3narUt8O1rvm++v7ChDl9WhokdOjiJY8oMxle9JYKfWpWkfsUPfQ5hmR/ohJB6pAOLo
YJcuapzCCP74Z+Dl4E72sPSHNhE72HBMaGJnd550H4623wcZlg1KnL3q47YSY3B1c0C7137kUNfW
lciaQ/P+GREIL80qcSm4n7kcFMgFTjhFjDiVvPLBmxyy3VeCeeSKhOIfvdA+WrDWnVdQennlk/Ru
YKn+2SdeH8d0eEzMPjMeqLJHVBX735jVLauhuLgq2hjHg57nwwOb2oOl7LgdRg9xwDWNxLgG59aq
ceqUAKQWFdhhPGAzApW17kFfZIaXqMihOMMsMwIeEI7Kjv7i1rBEMFHWIEyex47gvYs82HLJDerF
gDN6zNywQYW4tlA5cgggNu5YbsrxLdmGiNp82bn+bgcZZSu3PjFV52Wg7/7IIMjq4fDmI/2fythe
lyCVpg6iol1KGcKfNduI7pIgTqb9dz/il2qdI9jNQl8dZzVHrVCsAX34aVMp0edKobBIwk9wLMrR
3Mkm7rXTTXw2x7UOg1OUVRIE0AsKyPQL72PM1ybYJvBzLaCmzKAkJCs0Kn2XA9SmvwDiI6yt7+GU
jJilsEXaaAq1zWLxwYS3rLj0AoJRoKHB0+ny3MXtZnSk4gaLfYFOBgo4b7VIopX4aauRgDUkfQJS
LwhR95tx6G6a1j/WqNiwVPnQri8JjaAaXJPYXCI7QLBOg+B9FCcl8vpprIgvMHb0SkbXkw4BQCu7
VwjyFvPqwS70rUY25Zmy6cMhKTQzlNZzi3toGuVG75K0IUQNZeYctq5KxDxnFuIZ59Z4jkAB3FY3
7PweYMReUj8A7zuo/NHeGNwiJGcp1JgoUN//DOEjFa2cYGNg1X5rlzvObKDOX5ZAIiabDcdM/Bx2
ZiF8OVPL9fYUZmNOt5UA0oRd4EmOK8Vp8uLAe44GXeXmmd0dZH34eo7KoUOpY8eSBUcdAbeYZtE1
niILQTCmXx1CcGoyEpX1kfCLQh0lplzXXm5+ZLRLfCkaQVsg3rvzz6Pivm+pRIrVyFN5LBeOT05E
YHVBcxaw8mqyjhk4rVkCzQXKk6snXrYXSrxaMYNAVuwmi+L8YCBC9NbsSkLnJKVqcKLuEHRrFy6w
AAEgyYBtPa2czctlbpMRFj5ozfwN0Q53PdR/vlOqUzfYDf7h+tUs72dYHpnpHqgS42323Y1PjP5+
7Z0LRsv1TMG81VVSc6p2V/QjPmmvZP4KzwCCaO6xUL17PnNcnOeS+1RKbOeOKpvvsLey62IL/BCM
EHmZCd5nMERqTW0kp3tiXxpkLwr5OcFV4VKC4G/qP8YLB2fY5G5zm5XXuoyiytObnROjRpcKq+ue
abGTZBn9HpDwL8WXxz67i8fPPbNOGapesVlT6Gx2YN6ONbRg1SzEYzKcy+cjAwZwUHMDBD3fO4L5
i2KeDLW+Z++J2j+YbSL+KbJ+9YY4Hh5Ye8QLMzorzsbg1dwuS0P9wpveigJ9V5ngiSAXh4xwdwnk
gLyMcj5LJYIliH5xczs6m6C+UbihaPFk/jWo7lzDBnWupiRpquFD6NifWKkumRygbA8KtzXqpKfa
5aADrFN/jd/+geiNjPSgxrUkDQ4eTdibMLmoaWINyPCtxbH5R9wuSpCkxr8ZnJg2P0P2qrnz+Phk
3Hj/DH7W4t2N07AtjpxsxVKaMHOvq+Ye9DcQRiLzH9Cyzgpsylr8j+kkIGnI0pbEtC/QXqmls3LG
pSbwp3mtZ+azX93+dFq5o2QoqJGFto8e4JUdxw9O9rzkWeQ26csyLuuAGC3jTMJIG9s3tWYluDaF
APyBHYZa115MCzsL0gzb+QEnocgA793B2FknMfMUL5ZrcUHBc8gK+LOjgO9xV6V5cldL+ljkEnyn
g96WzGy8vfreBylNssMUJAzBCVI1H6PwQim3GTXvgW5ReZScVMEs6TIFGexhn+Fvn8SjRZAp1y+O
lrlsjCnE5HMzDcAFxD4hqxcxJAg2U87aEL3kuqX2i3uQHmhEh0RMGLnYLuccMJasXPKDNCa6urUa
JoShR0D7BA1G4bQl2O3aWktPFcQfQnT3sBiI/tNwSFCKFlNdcIYzZtpnYGGoVTyoHfA1i2fZhPPZ
L9YUwwjLYrjC6c6NBOMwCA1t0CjgalcI8syifABKA21ANIa/l7PG0q97y6Tiob/UEvbkXDakta77
XtaLxos2xMk7P8mefo7YmcU7kEUdzubtKQYyAX1ObpdMIdCRX+bBiCRjaPdOtibdVKVdEeNVpDQk
jtAUGH8NaHsX0kBz1Y35EPLna+EBCXYVSplkELUTpiSFXEVPxAlrunlAE7vMEkKloQLB6ASvilfj
8tMQ3XXSmY1nOpqlAHVk4/aOk2Goqkp9Zmseo1XnHhQAjGa6raAPHe67fMERiP9K4xD7tkkIBFCo
SI7BHe7z/utBB+prGY4o4L/71aroqCcyjQmLXcf+twywNkcsvRLTytv9F311VYMswh4g/KLZ3S5y
p+MK+eLglK07Ol/ckCqqx8ux8kDVyBlgrNSYxUS0nVkDlBExs1U5xRzUuVlPpz4qxnwQaOSgIDYC
nKpWdmabpbRrZALD77qwXEaugWUnf8z5uA960l8t5tkQpKXC9L1Xx6QcfOU7N1hAGUNQphw50tLk
h9aRb7Ju0VbQ1FIXpeesWRCPdGC1+e8l6R+V2PMY0tMDQ7aHpSCkR8VgbtuN5dlObQKpKvsj0R49
xixFgjpTots8mXeIHl/KsLrjHbyNmEoGHaCLj740zE0BcJCKCvlC2v0kM3B+qjyQPK3x1nbh5zXL
/yE+RbCpvJEU1TXi2dSLEdhe1fUIlWeVeE8AS54ISLLVFsFGhIaYgUxZX91sKTqG3k9I5FwIBpo3
gMD1ONd+Q0MqjqP978et0fWrkIytlzxDrcUwtXLtXRA1m8KERnerCGRtaa+8IiOdXBfXU3Y76JSY
5oKoffY8M/u86s9vU5cJsi6tjxkPZ0owSJfiVWwR2I3NfS1jcKeIoPYixZTz1PSdqYkUBHcaN2fT
/5C83jMRe4Y22copi3mrT4jKiMJbJ3velHHaoi6n36/o2V57Snk44XIbVUiqR7B6DVr/AUTj60II
T1qVxHYfUwGbBCkdPBfg2FtIwWWBxFxy7d/kwCFpMdmlSPfXo3gaAg18DnOfH1MGveM1ADxpSbqO
HAORvZ/3HwkLPJ120/EgsjlLnz81tjiGdwdvYyAbxILD8OXF9OTquSvaglgM2hVdAL5Td5D3vXsu
hxuxWJlCjKFgnbQDdODGp77BVek5rrmORt6NAZJljq3WmZXISwFMyIpPKlFfGqyLFI8kQgaouTuP
aVk12eI8UPrmey9/rRpxuiU9L2LPn8h2MilT8g4xTb8Db5jDfxhRDIepcqLdFjxr0QvsMWnUhnKE
1BJYU/yFuUlSEJM8+ElZJ6pyqKcv11jqozUJ6/lGXb2dWsmZ2alJ2qK4VSH9Q6hW28R2ax68T1F1
ivzod5tH/ituJhJDhWm/Llq9T7xKJW9P/tad0gR7fATzK4EWtqQYKj5lmp1bkmAIgOJ+MjDDAdIl
HGPjkGluVyl53yMTyGGjgJvSeWpeV0HypeiyK3Ql0RztaYTarI+K/xr11SvyZecPHGBF+G+2ngLt
zcrFiIWW/cYL5DfLh2Gse8SvPmXWLRdLCqpD/PBReZ+D+/lG5dBbSgQ4NMvac5CCIIEka9DwX/D5
iCdgxmOMCnfd4YwD9pV2HEqxvbz3QcxyTfcd4hm9pHhItdmgkZxFMLAag3ISQ/aU8EG9PtLzxmQL
kybJHTNpDqohPttKgFfkccjJ5sJg7HFAa9U9MdCxoytOrhA13o/Ay4YIMdLIdmneXH3xVaImmKLc
oNRVXSpptqCgDXHORE6DUcDdvFuxAyccJmqoX5FD0Ow7U98erpfIy0dFNpDQ4WN+XHrPRIBNfiLA
+VwM2qW8s0/SCfgVn5uOC8ajVEVmYR+KRZNUsttBx1cB2yApRakZ2mPNfKI0QERyL5GQUw/0hUGt
NNtDn7A+wsNPsyvPLvhV8/eMm3fOlR9YwxB7R221P0+alBUPdn9Cv+dkYQY17qTBxsgYu1NfWC7s
xHy1MI/OH9cS/NMK8SARLVi0a4LKAQGncRQnYrYN6XCvqg8jveLYv6468tc2eROBqtA4XV+JP7xW
G0frFgDx9wIAk7Y51jRtwS28CtwlhnNARWRSRy6m/9kn+n8hepqZPGTdBZSaQY60/uVinkdQ5yYe
TGn9UOPF3ejSAetpeUQk7fQgxJspXZ35IaitrNGy/9k2KBMRRsQIsT03/oW9nfYpqmNBw+BGU+4p
lZs3I9wj4yA6Z/TN3yd3Doz/FhYEaY7JSOhBbdvvAQ912eFW21HWhJ43xXjCgiNCblyzCS8xlCC7
R/Ko8ovoQTPEeyqfyEZacFhp3CXHcIP03yEcg35iKATTaVpab61sV/bOXFXOcJkJ20IWfNsGUuy1
wLgZO4BYFuHlah1FbSPt4/7nD0QKdt2bOmKghxJuvbE/cmXvjUyQsc1vZxnFetXcHSZ5sHcDkx94
Ckk44x0pcuyz3VW3esactJ/Vg+QoucwTIrHPofypCIGAwTEvH/s3/ABMAns9gBCDvxjsu5gSccP7
hjuNsRi+lKjw69sy9sdMSmVsk0W/iB20riwbPmcG/v1pgI65PwY6OLZ4G11XMRS2m4upxcUtvgeL
cSPukk481bTElJqgMoobxWo2TR2ChhUVaHcJoC+TzozOR3topsm3hx4zrniNwkz8NLCvtmRX1V27
+Gm3nExN2V0u22agv3ARDcgza3QqN6lxpDqxrHde8CvDat/jiOebm1EYePjeRGs30mS9GXjioStb
rLToUmsbfoEys9BcNa1n+IZf0kolVlRg8u1Ubrqo7+6zYtjdAQCQ/YVmwotsauD88Fxc1tNDQX1h
H/Gq5NSW3rQAdrpoCfsaxxGNHJ/U6hQRk0ErrJz7QBed2WhbTwM2qpXbOySQEAGXnRfERkM9gjAD
eA/JHOL+JcJH6rrRmKyFoBSD3AQBI/KP3cOZBVmSLZKiGdRWQDegD+Ocaqw3wEJ3vzSCNnTMRqKl
/f6LYV4p6EEqOJ15j80G9tk97THMK1krvsvPTyEeJ9/0PzeCSughwkdOOR5Zc0uISEhcBkvZrSwb
vx9F9ZKilY1ourLKDz9pLd3KvsFI+4m/hnT3ikNMeb9EJNSy6AA8cJKrUrNBPfPUo6jRaG9gkTDh
3bGnHv/YJZjqSkM+suY0dKYuAax5i6N+SgSH9CTPoa78awon54xDxLzmyOizHN1fW/lZFo5Dq4pj
zFt+bZChp5H2IRPAiOm2nGcELs1+IwEsg5SVJOtPamr0hDPAMmpp7H13AH/3asjf3yE/s4SXQILe
hdjkfg1ySt+IbVzJfhEl/J0a/r1RNqUY1k0JI4Qc+BEYxnFZ4UE7bw1zLHxCopESMxqI3P0iT2dG
5TssdbOsKTXaLRSSyfdXjZvrTi14+EEWYN2JJfT/nkR1JjBniMJniu7Z26EUq+Q5bDdcQU3DSPmG
0+nS3hy2EuCpqKlqvK5cbdqN4JPBBQMT2ky21pHqtiqbIKhj5cf8lOsp4EHxf6wUKac2X9kFOJZP
e/9iVMwdyjwgllzK8q9slkKjjyWJvGhx6zNwZieByV+Bv00pCPx5YxiYB0kSU6h8CUSFXrOJiszf
6JK7h3JpIJm6N8OHdar9gIZrD4WhxmUhMb1WTGs94nqDFsqJS1gh14kp4Kb7RdoiLNLRk7K77jNS
lpq6J9LOv4Q1GJAZrM9iyO9Cvuq3PshwB1rlnWkla/xUDcgZ9S1Y6opPRZS75PQ/LxOi6huhKEbQ
z8+pWunXVjORG8ie3EN5W+l/bP45/XnEceEC0XoJ2XgkOn+ryk4zYBsG4xsDiVQHbc2JnopP5diR
4vyB66X6yzt/zqURuYIfrFv4C9jHdta+PLsRpXqlbXS4SlZrhSeKqm1mMbXfaw/08tJdWj+ZBA5v
hWlIR1C6ELgxntTbuDgzljJgRHZS/yqoqd8KAw1uTGe9ZeyikOcOyAMhj/fjMB3c5P9bGO2WxsB4
vQiMPbxWZpp+WlVGxVH4PNS88w86Ne2WXOiryAyhxyO/SNGBKDuZMp+DQpOF7+vMzhjUrUjIezsZ
vLmbIJ2JDl51FNPbC1sLgNXAKug22qhRC6jfXgcOWB2l++4mdFW8Wiujc0rcvyADqAoYNlohWTW/
rcvWSIoAuvXKq0fCfS92Qu+mCb66IntesNi/BobfFzI+ncet6hS+nCyQqrj1FMxWF55mNp9KKMmm
q1jEtZN4NeS4QSZn/gMVtALrFqfOfkEMnntogNM4zyDxt0A/0I5kYRvlnY1NOmSRu0LE2IewREU4
ASLokrPA46NC9v7PbZNcryClXJbDfJE7OFMHP9ikvMNVlVzXx2YsMIzAKRiA6/0YvSi0F6E5H9RJ
atP1gnqF2jo/srcE+jqTs6qenIZJqPdFVU6WW5MJ6L1Fln3eHCE0Y5zPHnYUXQ0OQYFEq1CAyeSC
4pbgU60psSTCDfkvFYHBzVLZGe9bU24pfv7xctjh3a9WXQFFWPX4bcKe6ux94Y6Wpc3xCjT0CpWs
opmRrJnagTMKnxRSEd0DtDRvRFSQHepDqyRjb7FOPBWX+wwmnfO4cvBgGbzy/8YesR6gbbDNKw3H
b7XqzES41CtW8RuyDrol1pV4vKYlL/ukO+J2voU1fI/VoDul7YhGuDDysaqg1cEoiNzXa5pzrNER
lTW7ICsGN7OjJBvoqZTxe9sInBY/s7GoM0s/m1fpQRSixm0dslJXrh8RuEkxD2Ro18qH0RmzwWt7
MMRRk2jaCMQTFiJzmecRtUd/84r0TiBUVROSd8HtU9tnlt9PzTmiFr8OHFP6k6z4e8/Te9gkKCX0
MsnPRYrkVoLgdpoBsghA9OOJ+yzsfQfKJjh/Mwljj7m64TqC6BNmK+n+S+xZT7ml6nZk3rc989kB
PZsfGgJAWcO1FjIconBauiJBjC49qjeAkzztAzNgk3ptMekl5pb9Ut6fonZ/eLXLXqAaFUXiuyMq
jFp1rscG5MAFLj/kVRfg69QI6NE2zEvSMb2nLpljQC/CCiSgfKK4csI742cSKQEE0ko4Dx7k0QZW
DJXDmF8ov6K8WhjbCjtYmMJjQuFAUpeKP/tDi9O8aFWtNPth9tr7/ACAyvrte2PmPE0EVmnkmv2s
0bDEyS1SBMWPoNHNth/54YjuYRx/MuiI3kAd8oTyPxb7gVG8D9BELKWLYaCpsb1f430iqylwW+Ou
bDuQEf6ah8Za1ZB3Tgh4WehUO6PFYKcDLpT35kuIZDC4TUEr/68K88PaqZAG/FIVBlekvSDWj/di
vlBDxxSuugA9mcmOyLSgUj3bHYPEMnlD6eSJQn9gJEwAbFDrqn5dfG1+epVKAqrbEIHiMVdstWmv
J0CL9z4Rft/aRq6hpYjfmcKix7r6EciOlFlG56zQ9bDyCwJw1CXf6boezGgrM8Rbgg6SsqZ1aoNX
DEO5EOoysqqX9BxbC+JNrxW+OZG0QasoSKrdLg1L3rCco+OS9aD9xING1j7ULs4nktG17G/uyqrp
TqGvwJWrXgknNtOZi2Rmr5k4xsjIWGy8qJbxWdLX7xnscQs6Mzc62xTH1D1bPhe+xQ54vjtJF9af
gL02U+mbIEtrE3jkgEW+9DOpuIFyk8/1OY+vnZn/vJ4ffJt2YCdHpyMN3hiqJ/6Xs/aPE6VHfUyG
00/oMuwImTBUUVbF6Wf7+mVtnZSR8coYE5vKErwHHdbW9s+1wjO4hQFVKxY2g4iRZuO5NkqW7SAO
eYOgg/GKtgvK9Yndz3Q5yD7UbU1vpfcWV2zGDanX2il+PH98uDmzdeIYgTrAj7L4DrVzurHkU83y
CK3b7zM6r6CFqh9SFFPubhfbNir27JCna00Tuh8hBvBNKtwsFOsAEbVuAiWyS1PydV0F2ZPM7k7G
Oomn3xFHJGDORCRioWVfkGedujx9g5Rl6VVXyuOdLoWG75/5rI7wsZWrO7xNerhnJnEPxU793ybS
xgd/qyet1eJ4KqwLxdcfqv6cyTknzWH5RcF56jth5xghxwUd4ov94hYFhLfOukDJ+81s1rQw/2vI
4U91m+uoyhdrnjZRfwDzdI/kAOB7KeCuyd4LWSn0Dv2f85wwYEZZSMCcyoqVEKV6tNWC5leDYime
uUVGHlz92t3lEt1pbni+TNgA/0C3ADoVv4k65YvTOOlhQmzVcYhHe9DcyZ7ubkbtTxswoN94VU9J
gilLhBt6Iosreb1el6Z7wUngT3s+sGnDtRZeWZYJ7EcRdp2aVVEEZc8shh6ZUIrjGUbynjp9JuZS
gIyFpTkfC9maz7U/BmbwwHZubwjOplvPFFJx8mEPMP3arn9PvKjSiwWuGVhLUq2B+rgpbJaRf6Kg
SDtXEZkBoB3vvWao/uAxLagX+55+gFVzgt8igC+XwNK8+Cpd3xTNjyzikurHUhYMf04zf+EKNd9s
CKb1RKxJz+5FRujHB/MPuyiD0kpTP0xdCxB41aEp8cHwxkNJOsfOqvMqm9XspaLVfFqv0QM8ti4/
cceOJ5ecOgAIEMsAlF6eTJmSTZlSNadtR3ae8/rBPAOCFHpqh3j+X8RbyBC1MCPXSGhNhmd8h03y
fN2rlDuA0BzSAh+HLc4K623lIlsN00hzDWlreDiPRzEURbWwgvweG53yQmw0wVpPJ2gRJPNrkCDH
595w4wxXgLtrpNp7JwoQBsteGbfg8P44vN+WcEUgldgfapVzIJ/bpGgQIwy40EonXXQqYZmle08Q
HumtMIRA8gf40Wp0skZ/EMbWDTDaeGTa/r1ePtE1TZLzZFJ3itPTjujaTlVLBsbNHvQCi+u9Yzft
ul1Z9wg68n8STQDUkEAPOqyNmkjsD6OAmPlXL80+KJ7EdvD91Jl1Uxi0OXy8ctWu60m9FKN99bpG
iX5B9dHcZS+EWn1QkQV+pNLbkpDy9jNThoZ2UTdQUbOQa1teWfzn7p7iLa2GbVoa8GCrIfRtSHdc
9fF0s4QSuIG5tES8ZtTPj4rQRom6hfzdBaGTffmQUT3a5mDtwtmqUKVFMq/IcBkYxN109Q9yHcPq
avSrHILorvvWKpPW/u/nimaCSslSeKq76mCgZP0wedSbDOoJneRMC/IijawMmjuZMySJD0Oxks+a
GeAJiLv90k35fGv7/AhFFgYjQjwYIf8Xb2iK1COmZ8GWX7zvEVhBLXemDEga8zKK8PEvyVdw6oNg
vWbbt4WXIQ3Kxc4Lk6IBL2JB7V6ymCS0ZMATrlKJWly6cuUQAWe+GnXPG4WNBdjy+zgBaw6p5OBk
9xDwcPRZqwD/IHKxqAIqeehxQJULfG9PyQYy2enUl/iWimmTUhYhDhfoqXDvzTET311Ek7y+MmKB
xiuHfKkfjsAISgp+oNIW2J0SYq9Nd1ykEWmhrGu/mcWW4UnciNxlIEHGE3yPYGfH2Rmwv+6oYQKv
dAHGuoglgidLr/I73jKWtab/zyZTg4exA/xfMsrLJVBZuCXm5Fi9Uy1fvtHA9YEzQXsfva3XY4O+
mSYMWcN4x7Q1Iplu1ig6ocxtElHDTJ9GoL7gqDckW1vepCC745msPh/wkVZIvWROjQVR5UoBZOGJ
m7BJEaZ2FlTHaitsABYLGMc/3BcQYfTofYwWMJRV789dkhFAgnp/9IWZIcVoYkL8V7xbkQOJYYFT
joCeS8lCuIEyGkTn3Ucw38TpB1e44bIzFcIv5wmKdreJq6MvQ3C7pJcJyFVyszih++ATGktizn5o
mYWm24zqqb6r0iF6kd3l5WRfh5dQGHuNUKN5GcXhDobhPOANMhPSgnjydBEZKXDzQtwKhqm0+0f8
vyX3JfzQdA0zUHZypfeQvAfEE1fTSgm0+4WhQNew7phC/D/pJFz94etXxcqdE9J//Bwou6PWAGDw
Ph+vnOt/fjutv0Aa8xu8MzYV352RIKf1FGVDDn8o2kcRVQ616/QBj7ab/KHkdtv9q51KVdskWjdX
l0igeAa8m/eOybVRD91aODL1cyM+3zSwqXcDlWRku5VvMwbaa5Ek+aWXjwcTKb3pBybvAiiCR9C4
A1sxD8SwHiKhNvRipN4BKxmpCeKjtsk9RKYLvqnwIDADMauXSlk0jSjAi2NEoSysjJxTb3gMBhLj
H2/a8WI4929Xggk520w1Vn/XTC+iGFKxZbDMvtrHbOzTkUxHxHhjQOFxPkT+gx0fj7scTk4lBUBh
WaGrzJFFprnWOYrlJ86YocsBRoCo7xt7JkVMZo//2WCsUmohRebqcP15Eskk8KynbxchGrj8vIS+
cad4DHymK7Bv0cUw72SwDKheJmUi+7i39IK1IZBTDMyXRBxdnJ7oOKcmcuyXQTLY8b0tsqHCd9g6
+gc0KTz4MyRSIkAcME3fj8Zjx3GOBGEPzWvoMS2ds0JJbAv1o8yZRKMdJSMiB7DUp/Rjdf1SaMLh
RkqSVemdUmTxqYNbFfYK10Ol6g4opZy4vRbRTDpfcPkSkgKLNDScBohErEAjQxzA9vCdq2bh52j0
bI+R1FwIRMO2O/dJo4X3KR+4e50lrsZEUkmvWaj35VeAfvFD3SbaDqTSJExpaw4Zed4Fc+3oIdze
yiITnq0dpnwjOtun9tDm9Y6I9aZhY80NrRz3+mjh7laihLCKaYznO1Ms2I5KMDPy6UxV75Es+2bV
hRc4gxmsAPmaqyJ65b1jW8/wvp1Bcyq/f/nj2T+GS8leC2aTAspZvFr7xLpfgEAQlZNhTIVASbGT
XzJIQpeF915VlmpsydkOLtuDa3u1bA3NSu6jZ6w6+GetikVr/KX3tCqxRdmJVLhEoGs/05082JP4
R6ts755QkVLC0kUjWsp61xCANf1DpRRmBRekLD7JwcElbUAQ4yzvUhYpUgsgh3Bg4dh/bHv3a9C6
aXgM/kPheR9k4T5aAm7c3l2MJ8yobjf4sXIMaf+nAmH7krr5kc01fGNzvAJELFGezhEN1UPGHdS5
STdZxbbQpbVc3j07sXNH7l8mHRd/zhVtvqfP5bp363XVtXrQ2JGEA9u2HdOD7s7a2TK9EwicHWph
ClWRxaehdYKGF3/YlcB+Uhyi3uDZevVeS7iQwsQu40Kraa5Q5oM/JmxIpnmco+Ww/kv77OL4rgEu
e90rjHPICICnrxVxJXCrsMXL9Qh2ZehYHps/ikenbCMeJZLlmbtkjjFoq1tkflHw1MA17vamNxyA
R6+wo+ea36R4J/o/UG2j7E6UL/JDtML3CLD2sKMivPbCBfeXeCK5KujHZozzWvAcoGUty1jPOW8V
nVc1Ac2I1ocWGlj4VaKHa61wZ9swhxhP2nGHWLbFxZJ3wlGVTNtzl4Mayc7UKMt/I71Hb2YDwMZ8
XH7wIr/KiHKYlekFKg1OGVaPVh0I/fOJ+4ix8Usr/mnag56eVGyjpSkrexdXX4IfgbL21gdrj8JT
3LV9Eqa7zb9lNI/4K5dX3fLwa+M+1jNc0PlEvb6pb8YtsxgRfi+C4d+NVV+YBwJPjTwp5JIfETu/
PDXgww4vqX4SyqPVgRybsfiw3b0JwOTgHmlQycKR8jH2+nzYPeDBrSgMg297uIDjWfYRlgzWLlrT
SXc7eFuTlABHGG709O5g9KV3T1ouiL8z1jW4TPaYyL8QllIu3aM2zsWifNA/lA967yg2V8X4XU2y
0A5KirpW6j2YFwbnN9nXMZa1RaUMzqsbeZzdRLCeb3mK6DyHkFtN9V/rVH1MTZXPIUe9L0MoDm9z
KKr7lvuJsGvgTopgeLzTLrbC4uHZoVff9bEuMsTu/U/K6H6ix+EbFzojF+t1fGvqNqn7rBfAtfXb
mC2X5hypS3LG0a8dZAlSEATdCZACtKEGjYzeuByUQbYHPquWSdfms3NXudKCLp8ZEcZl2ECeVvvd
m/M0lbFpnX3DAzF5i1zCY/F+9+8H6Q3SvHiPCVZpzrbfSdR9O6oHGSsiG/1xU4jsaYOhdV71QEWT
TiLE9xDLJYwl5lw0ts26YUszW7qhIuyw/JTGfFEOd3VUxtv0Mus+IJuGdHZAnGZRVevSjAd58klV
NigmxunRB1++3TaUsz6IDt2I4DOIuiCMUX/TYYeEG2CD7vlxhcgoSG/lHLZWNTluAIOixuEe1Sey
YLSGChknmgA6UNrax4saTc2DWtAAybGsijtldMxLU2i6/JFvZ2KBng08CxsKzeQkoEVO/ifEDqcZ
YtbVTKQ/ZH7dsV0FYiUUOSvu/45CGcpyssE5VWRFdCYGgffJVF2YbGiWGph6UnwOwqkAFflaX4Al
VcSdMGvo2OFyMWALAp3pSQ0FuijwD1skqP3xN4lPCPYo5lycTs09KMaHnoiX2rR8rI2zEHxDQfb5
MPf5aSTdVAAwPBjk+9/Y9CHdV8QMuT1pJ2nl1U2LR28bOGMOH7N1b74mtlN0u2e+N4BO6ddFWq9e
x1TmPo6LpYzrHYVWHbCblz0DQd5AWBPVVzK2TLa3OF1rmTN8BsmjQ1HeIo1qMwBE9GE6TFPzTA5g
IvHBDVr5lHWmT/05YuaIe7RlJJIxXndZ2IB6E2r+rTY+lMY+YsEl/gHTc/qz+/+nlR3JgiLsnBQn
/Z0atZK3Omzg2sCYwB1Na9YcCAYECqSGiT9sanNUSO+6A+ua2Otr1B1MTmf9p+03R28xH4fN9lJl
1bP2grWyQf4B9eNE1O29hov7N3t3+wcY+6kKmgZYeymj4ij9qEUsHmVav+lPC3mYdBHghF37Z6TI
xauM3T5rtKHQFw1jDN24b+E3UUzjGkujMQHo7WfNDXHDN7v4uGtzTUU8OrUy92QWx2U096E2ihry
wBrgJQYWGyc0CP/kOSj3Q1Dw8Wr8Z79rNKx5MYB1EMG3f4i3K9Clv2FLAPY+0vXKu6cd1zOtM96D
6teOOQyzdyOis/Cm9eCt87Gh3s7u87m49E0gJtMzwkphthyDJj8J7DIqcSHouLI6QPUPi/YZfkSq
mZsylke8+kLNo5Ro0zJDH4a9sgp9CkASZmLui+lOQwZkT08K+kzvPfRsp8oPM8CXcnL8AOENe8ii
CoNvrIi3/L7sz8YryUCxayaE8gM/2pxvOJus1QHQ2bYkDsCU1mXWt2K8+dl1CiPM34IKYyBHOBNx
Wf6hJw+AamjZo5YqsnrKspwR1u/Ldjw2SmflzNxrNhaCxvolhEqIj+dNDrab8uVDRAv7zDdnSWbU
wj4li6r7sDFLyhFPymENJ4vwIOMeJAmKdeOd6RnwHtEeG6O0OFjXRKcI/50onNsHqyaEeYanTz5D
kSjcQaajopzjwEMl30j5KT/pUIVTsJLzyLQfNer07cHiX7BQ2X4vyE0kmhT9JMzfRSEbaGa9+W1C
/rqUCUs+fP+NshlCbAXfp9BBDfF9HSV6aZNDLQk44vgzS7CQBDhg/MWFh18pnqKYhbNs6sOzCmUe
wDQ91taKKY1yHx/Cam9XQpja1xlw75qDfFFUW8qNoXMewwV9OQ877u9i57GfVJxjZ9YQrlvF8bwy
u3ag7qN50QV1GH/g9lGDLb6zhYK+3mnWzE/d9CzMjssxPgsosGeprKrRcDaLA2rptjMF+At07tWG
c/VKGJsVC9//6ncaufZGpw7rJtiMZ+fZBxZguj1LsLA47P/bfVk4BPKdxyDpPFaf0/9Mhl8qt9cK
Jg/sHvWwF0N0/jZIs45wo2lu5T+SefhvpYpbJmstCONaO+ea2Llk9DWUyWaoTFR1eJA0SYFTG2ga
hirLu+NIRa9q/I9gNdIYq7DqWt3t6oeuNpnhadWj5pRAE2Qad8EwNKvfN+uluUpwMIRfHArY+F3x
zfs/jL686ihrqwyp55F7OevBRv5CI8l1zyEDqLLXt+F7voeXyEug4ZGemF+N6cpCN0AkwHUju44U
1i3VK+hDhmLUMZDlUNORKu6d04GKqKrZC6+bSdjTaguEzlQPzVjlz+sNlfHnzHcAZNsIwtmkRU8c
JZ/Wan/DoTbHN293owRc/dwS/LsDqLLtNFphkb7hE8VpkhtYJJ3FTQwpFCy+MEow87dsbxja81WE
FwkO0GAXDO8BMXZrIaVrloOvJcshSpYZFYQd5KnC+tDV04aPVR23m2zYBd143nOuUANg3E7gezJf
5hVC/osa+cqERhK2Z6ZdSYD5tqCZMTxxE1U41/bHnbsTIECrdkRYnB3j7W+QJcHfnAf8HFPyeBrQ
YApBTPkS/d6HmVpDHcuosNFXV7SS0NMtSLY5cAKjEUGSX5qP+fQXCOILG3Ua63TLxZPSckv0rUHu
1kaNvYT4jh24AT9C34n9d1tlN7B3roe0ETyIa0xmuuhFR3YjzRsys4CunTVaEGNCjdWMWW4mEvS+
LTKqZebRI6IwHJAC7x4OlBvY4fqxcVGM4SLKxDPz4f7fOBfU3tg9/3yCVS2UsZB8SyL4dTIsqkyA
aojbv2/kMUdHgnAgaAL4DW5wZ6jpTOkJ/8I0Cica9JQ4x+7yTFV9/yz9biFpJU6+GuRxT5g3K9za
+Bak+d1JjxgdyIMUqWylsb0tciCQgk1ur20pbk9OkkAfJMHEZEuku3ZLQaD+hm0B3Xel4Z1LxyC5
4/8e35cqDWG/W6xYiyMOv0LwnCCrDZviUoduDXv4t+nqYn3YHhdKd+gdvMDJ3ZbKgFeHz5rQNWjc
uutxCLhiideo150pCpl8Jw7s73Ac0ENTm9+QB1VOF0u6ANofeqC3z2xUr9h3KK/QctZU5+aScBuZ
4PTnhkn5HPToAuK0fYNEFEOTLI7b2O1Mff9NZ85g8EUzseVg3pkADaoZFLIWQQbo2w8fqIKKRet4
vBNwvlN0CVItpFmPP3cfZoSJxPO7iHdQKRQif6FH9/aoU+ADLjev1hKGh8q2lyAUdT95J41edz1+
yP08MHopUAzY1G2F64Y0yS07hwBIRLNTDJcbatZMpQddiNbsi77/NfuPCH6Pr/yuMN7aAUDxAAJM
l4sODGEPsdhQE/8pBF4MejXNjILuvuv7wLQNzpF6qKcETRXSd0mewfVRqkCr2gpR3zf7vjHxosE2
k+qWs3GqqmCOM656AToCSU2S2t5z+5Jespfu8cq+ijyYExtmdTfRaJ4Fg8CPaN2BW4X4g2df2FXF
onQy0v3cYu3Zspqq5BOAtPDSS5RQHBLsT6RVqxoOVyX7vnC8B6lpg5Jam4P0EnxWD4yfdKxiVyaY
iGMwnF5a2eNE63PHgnXUDbOnELHk6qi09Eo4G3Pdwh6ttQSFsOcsigpWFv0lIrKYYOTv8JWnYEfT
mpvS08rgofWEMRD2hj/RAheehk3oUXOcZW7YB8H2ZIZKgbsQiN9ie85xwXXpES0PLaShaFWA5J9m
rT47F90K+L0bFP2UrvXlxv32Ca9WKQs007cx5YGCSRZSJueLTrc41igeWtz5BQDJHHS65jULPIzo
Og5TQpGtGvb5E3xiYl1PfXPnxoxg/I2Nchm8mDqMD86IHrONiIG6BrIakh1Vj0KjXOgJQusDUOXD
hSUr6HZ5BZazvF9aH0LYedxSQPhgLiLvlqNT9clDiwHs433r9DJWRpoehnAwpWGhGpHwIjlpu9FK
VSM246DtPJll8E8KUVxdzXz4p0cgvf7Vt1ZBZvVSi/snRQ/dCJp9coprvzMnGA61Y4R8IqTugl3H
9cf6RvjFXHxB7+CM+Yyc+vbPtLzW0uprLmo0BsnDVKHxspj+DZQ7ku1LAINhKCrBzmxwx4R9tPil
na4JZbSBbFsyOF+ATfzPNY+5tbVEee1ukSPez18xG61SwtQ39VP0F2ei2+8EiSGq3rWb9PmXV1Iz
XLfTD94xw/6iJI6/Ayd9OH/1hwuQ9NkjqDf8GlW6IKDHpOWoX7D5SFlS0D7pDOJhE9SF0fwCcu20
BiDnKMxmzmzJxwNaUVL0awkU1Rri0qG2FEIcVPgbhVT6/WwViBnMPsW057xn4Um16SVgBDYACETU
azwNRlDgxMP/lIzdUQYxYTFaQbJQ8N+BBMBftRWOuWBsgoy6mmRiZPK4q+jhvmnyUSBY7+WPTDZ2
bkHNxjSBJIXANE9Nl72XaA8kKVs+bAs0sADaBMGbCr+IKFRkFAQDcAzlImkfUKegCI9mbPRX5/Gq
8dkP4KsBQPak9VXA4tRGQeAEDH1Yc7igURmGRKhY9qX/Ynw97s1GixD+Y9WtI06zw10OXWjivI77
oDYzVIpsUky6UqlUyKOCrfWmPtwhrRBXY+BK1w6qpWMXieIDQeMyisBoULp7zDVkCs2aEMfgoluH
+0GAGpJotKSuHUVWRID7z4zSHcTDiV+54x19s9FxSSONOymSONtI6wN3npR4vwqfGOlzeJUDtdum
PNJSu4V/g29lanajDEwC/l/Gs+zqaZW69Ntg9T8+5U/ubmhP5aydA+ABq2eEnxWZ8tx+HQx4nY2S
2+j3VvuN8/xiFr/J/UZ1S35QTO1vw0aJlAcmWfbNiFGsdAlRrnxylUDMHZveKI/mttLvFZiBxa27
xvpxSL0FpvJqrCXtVnMVxFUSgo8lzFd6ebZQ5nQ5PedCb/pQDKjSTGPjuPYAGsHv5/VJRGL879bX
COJP5n4nl/k/Zl2lnxwIA1lIUi8CWZn0EV1HNF1aXmIjHQlk2elD+wG1gnxez7O01YM9Sx11vlF0
9v0tNFQvjNeYJFpg8WI2no42LZ8oBdEhc144kyAR/7QucJzGoCkYbNRhI9M2V5zsXMIThuEJLApe
Wiw+rQkBr6XnZWj6u+mTUhMgKJdWSyAP7bylW0/Rv60k5LWPNk4MCbfFbQemb/qbwrrsaLusrI/p
+kiLw+8CHvdA9mIATbb4Q1bKGvPHmUsVGyS+da1UlmpXOzjXsf2LPQhM8WgHFo/zNmAetnQf/53E
6JKIYXdxa2iDreqUbAbVLckoVhBNdiPC1UxV8VxZmprSDVv9bXN7wzGWd/fq5On3WY3YHGyZSQuc
yY0i7ZCqhPyB/UQcKkZWJ062TTOqdVJFhlnQBtEK4wvrCKoOksWonFO71la82/uGXvjpvWReJbCS
MojQbWCOE2chXPof+mRCF/JuLFjfYVV0Wfbjhyvso8yFwIyOPjMN1o3H2fPA2jgeJyrLMZ8//25O
gqLRA6KM1Hw/tbwHiGUFGdk1zGx9YiUGjGPJmUYiCH3fu5KeaBTYnDq03yMSBgubYL8yN8UIPqEM
Ntwtm4+yAA0vy6oapWY3gg4OX52F/JXD9LWXoutCSQq9p6FGZTaAgpbQPcmTVHGkXqYeZVwMP7Np
+BO0d0JAym7QNktC1uTU3xOabJXFIm2Yt7zkkRzQ9a54jkojUGVE/xcTIv/DyWkCt28djca/DbSZ
lLrt537TqLCCYBvs2xP8w4FEcvje05+efVwwUn9G9xH1JZCUNH+sj7ovUvNGFcAupniS/j3nJ8RO
X4D5yUmbOH6r29BKyTxN97kPHUdoXzzH+j9MtwoEAzympNDGfgNOXpYW6oEc5rvUNMCFguasFhXX
279xgSntU43pFOI3TgDeX54j1X+b4dR/H7Yx5wbgG0iB9EKhxkwzU9XvhwrMYVa9udQ3pLF/RE7M
5huXfdTmSvC1X1khAdP/80awp3AcHErwobR4WUWCN1PniVlgcs4H5SBsi+Z1ZDWqM5qD9R7VBrVF
7y3yysO08kUoKJ83qLcrMZhY+jaUli941Nq1QHDUu+MigVCzT8E54z2gN3fY5bjkicCtgnsNSZD0
0nkKLa6DGa7SxIce7NV7jnvCnUiGN/wCZryKPOFjF6oAqB+fxcQTYvykfx3o7MOKdZjm0eK6UJue
vfxzxPL81d/0lZQKucriEacVZc7P+Mhcg33t8f0xfxBH+Ekz3YTFaqtq3Psblf3OKnolCV1BrEhn
Ld0cgUQJOAtl61Ilx3L2tXkpCJ8eygO3mpjbGnvSN3Y7HZpCIbCwXm0zq7tF/x0xGjNUITe/yPfc
GuCtf9s0S7c2bVHmQ0CwMRY714TbOX1xF6OY4Dh1rCF3/N9xvsBfx7oAsovkVAUJJbfkJMh6sA4p
P8QN+u6sYDQHC36px8PamRCnZ2sET2TKe83hRL3wCjtZAbRfQUQoQiFjvVdAe60e4iNmXe7MVQju
vKaFmKsuQ+14QUWFoDbn1hLKPZ/0Yyb+WgHwPa0+gL4QWdhmblS2S0on2tx5xc+/0S7EhU6SA0BO
gcDV9RgDAu8El6HUJ3ottJDpV1n65pFY9gq1fwGBH2d6aKMgOg+GXE0BIriNlptb4alqFwBkKZJ8
ObV067CrZ4YOUBObO3uerGW7srZdzH/LjEWZ9vUAvT/SqRoLIm8+w0wOBFAnrdlfvBBYyjqAsmf8
MIxlwJLlApDe/84pJnmxldXakzJhA1wkfTm5UlclCrSzkyIp5XIqhEOhpq8BeI6qsjM3KTpRkVpn
hXbZ6t5EEiPnxAZ+TO5OTpyHCoCSSP2bncgk3KDUY5CO4m/SgLPW88e3MuWikecIEpPxMAEAOIX/
RCJTl5Ao/xpyl3E3Fk5quomN7UOKIM1yMuSaDovsqjz4kxXy714Gk3Ts+3AuD6COwvQaZdp/Ivw7
H7mD5dRIyW1er1ZF5tewsGa1VPiZP8VlEPMYSRS1Xei5K7wRzkvcgOx3yS95bnuPHnotNDzocplv
2F/SoJwGCgQhP4p1jP9NcrtllW/I28jPp4HTKD0NaxHQQW6ML5lFJW/OVKYJyfLil8UBY+qp58hI
CBBDq44y9OYqAvtbNIo7W/wACHKfYp7Q4YLXHQDSGYhT8dfC8fdtxKpPH8rUVKFXQOHw30idED4S
paL8Ps57JOpo9NUzbvzPMdB6lQcAQtxWllfG7x7/Bqot3TndOnbTVnCypY35UQ68OqWa6fGaByyM
Hiaf4iKNovbuylHNXPU/fcsh3GZWINSiGaa7DvW7W2qKL7mHCkhbFsYjizsSFCf4zHqo+lkmohsW
yN16FtmmeFSJj0nRKg2+SreEcrQm8ZCUwYPPGSMk8hWhC5hxb1ElGDQ6pS+spDP7XpKYmpMQ3m0u
XWfbyiO512mM8+K3r993guKBGv9P2WCJrxredPzOEToE5zinOmLEHzpqaT1pUDx/AxUk7N5fCuHz
ef3RxtFD7rQfwwZOm5RATKA8xxXCQd1/11zXDdicc0PwvGEoNPmzj7MiIlIZajJdhNCRO7Oqn5D7
cHB6eQkE6SL/WLPcMr1xqgKaRk95YEdHIlHxkiWuGwaDKD2oh/AQUejYLwiFv4B2JFKb5tdTjrMI
IC82770YAJJTgrwAE+h8SSrZcdBn8c2RfgVXcpmByMJq1AQF7vEbxNk3SzaapHCq6IBV7rlCO/aT
FXD1ArJ2BvtLCG61WeusG+JL+tXkoJtAAeq0o6G6PGEvOcgWA6+h09jNBdaLPSql8UEMOzRfZzXh
0NrYA7PhWMs/3nMC4cjgF/NTCqzYSfHDGsfcAhC3AOt2Sc71tUP6J9HThgsL2Ma27Lkwd5tBva1Y
xMHMTIF7FLZj36i2L59gIdlqeOD4qL7RnImTLtlWuc1Oag3rs8e6pFxLdN1MK+sjM/mnn+ryEibk
fZsds5mC+xoVAAql7EQExe7ijlJvV8avlETFFx5puWchDu3kWw/DbVpECpU6L3ytw8aGdzmS21yg
u7rIYElwasZcYY9r69s/VT3L5TPxAfhTjrEtHzxOM6U5yc2stoPxP5hUBvVVSS6zZsGLcQPDUx0R
0OgP/A7q/2yS48HnWqEwaDndZz2TMjIxYS0AtJf16ZuawsP4Zbu58Uh2xgghaag9GBIQm7n9no8J
BNTfpLJgdOvh99Hat9Nw6thpEMKWo+dwy12zd8G07xJGexcc+zw1Sk7wO5cApXph1Q+ZgyJkfiLb
mAdifSH2tUTr9o3mG2G9uxpe7p3OLESm7yxjDqwDKxd97nX1TNB4GuVTPORcztp2aF+NQx/Szwun
aQQ5HRhfRI6FOLLHJRSxjtmFGNpHJ+IYi+H6qBcLtSRnp0jICgks7h6FDFj/trcFqUtBUCLaADxu
0mEatZ9vDABZBgHFp4o5wKnrGYxdJdtirpOqOAbDkVBg0zPfLSatR98/jcDfGwywF03rWcZevxBm
60LmrAWrPtQO8hC7F5+Tsir0PFZPWOKOVeasZwuvZ4fZB9QBVeGDlm73w5vJS0X41RLSqp+R39Vj
uB3h9tTF7iQG4liNB0WGkZruAIwgaMdvG1cN86bWUxuqQ5Ii9RXJ3L602dHodSSXWrEVPcrIiaNp
MEzi3nR9rfEJ82jquHvAFUIzJSVoy3xf9V6sWYuOYgrP0oaVsLwx7NV0/ERE6pszov5KHEKZHpZh
15XHNts+5LcMWnYXvhPHqfyTEmnwcZTSs86NHzTpzsQQnU9eqCArIgf3SGhR17jc9ILZK9jC+jqV
Hh25kx9iVa30r3S6j+7cPr62YMFpG6OB4e6TyZxGfF/HnmzwqhhwL0Z3zqK0ydPBnhABwN6+xZhR
8JjUY3s0icGNcoCBzn2gxKyzMl2GHcZ+8Cq9JlRKZrmZn7PFWyQb0aUShAI2IjFPB7r2aglOs1H1
36gR6HSY2E3QK+uPYBDAcTiS2I+Z1GvG0Khzb8Fz0CH93TSBj0cECpR732jwxEURMIYD1stVTm4t
+OZvo7GCtNMmcEap/eVGMxwlMexc/41eiDMYRZfeOYL2z3PND841tO+tJ6sAGMzUkgJemm1k2MnA
oAYZktOxGvGIsk/a9Gmkxq7sE5X/G2nM87eB6HvtcL2DjlsPTNdxMwwr1fseackcPa8x1bvsKGol
SRf30zklGpnlV5Gxs/UhIPZ2BwSEnnsuHJVvGVRWD1y3WleR2w6FvO/ncUeyv1thLet/4eKl4UMO
gL8LWXLokhmr4zXEExPVzFHpsbZ4g5U1V/rsHGjpiD5p2+okI25AD2ELedVkodGNHKbL5z0H4zAX
hmqmAayoOA3cIACA8/BPRmVkSh7e9QhKp7sSiPFbCSnTDToT1rbVVfKvVD22ZbDeN/f8HObdPi+C
Z/TN5ReZTgWFt44jFOrHLWJP1L/jO9p/Mewftp3KZAbMorf2sGEi4vzbr68sbd7qZ6h0ZyjtOMdC
hiKj8DG+KyR7M5ywUXctwElZo/t51hGFnVXxRg+8YKaSTMW/prHVJWgJpCWMNQ7UO7YiTv8U+LjO
9TcsA9rCvGkYvdqL3i64h7YsDKBwCNbMzihxKJ3xzCyhoErHd4mH/OkQNYaZEt2sAEpz/NidDQEF
QQam0rz7wShJNbv4xW5JXccPMlYBIkoGJiwKeNJ4MSpgjIT+kryacV3WFSnqoc2Ic6BXNFiG1W9e
IHPyAOLBw8XKz7DaLCmGKQ+0WHUbAvIjC8Iuf//mn+u3KVkrhVjh2yPNatHJUqpdACHCAVzKcNps
OrJaoA1O5u2SMldqZTrVVyspsIhONFJvXPjyh7QaJj2vT7kKjeGIx57b+NYvHylH1h8WgfAWqcZS
JlwtDvOeMwyeomgvsiOSxcbKp6EMPotNMbK65MNXqaOxnqpdOcot/zEtTd5ePFXe1TfKSNDtYaNA
vwa43QPpFcLbFA9N3lLdvpXgA20yj5DNlh+g4S4RgCaubBPdDdcDAUFZaU/LQ4O92pJAqUOO/w7s
s9P58bfji4faFjbvbWLOv5jlJWsM4zmf18aReEJehSn19rofH/YJAIFZ2RRFhpA/G4ViM4tl25e/
+5fTvrhvoTAcqfGSi9c+dr9N7qokdy2u48EQRuu73+mtrLrXssD/8heW/RwWfld7FjI/HtmjlUVJ
NuCOUrX1seDx8LAJXVkkTSpJuSiEFc80CMINsiab1W3YdD4q7yiu3LuX2NzJY2X3jwjC8Wh7YQtX
FvJvuF8JM7t8x5E+/bHPB7+dkpypA9Z3EUzZHiGaNWlz4MuFqvPV6uoennsHfGp/FNUzBrDf1Cu1
9ePych93PfaeLCkg+t4EX0F68tdsRFsc1Z3fClgIYiPgmzaaP/tM+eaXZhta79H9EaNB+iPLJgnb
Sj20KmF++Rlomrl2fV5b9QQlDtfMP00MRMuvWoszXgUzSTtY57mi06dIEaTMKfUcSMQ1HFwwAwlj
HVR+8aN/67+JB5vwb20/6s4KNkckloT48IoYHPnVrWQF5ADZQ7Z1CUoKR5XJHPOpwbAMtuMkPtPx
hXjUF8X+HkW5l6Far6TSKZvXoRGCyHwtxeHNDUaRZaZOBHp+qhdnCq0bU4K/H107vEK6l0bHUTwe
cWdRZBv6tZxBf64lXkDk+o/HX4Ss0+r70nw6f3KdcrDtc1xpi1DoXeqCF8Z1nTiud0Ws4w4FJxVW
u2wSDzWlOhslkOdFExlCgI8CkLU++UYk3eHcXqZhNJR1AyOal5rzMv3FSoeCZ58/q2Wsp45s5obt
RTieu9u/KisoxYfAAC8TjH3ToVcf5jhuJCUR+ceUcny9OT/dOObujBB1G2MyYD1lH2EyZsMjaiXj
Qe54E/4zvvUbGokAk172dc7Dl+e7CqQTkILV8dSaqsaxU5zoQ+S2411N7cA74B9CE/WFBQ+wR/AH
9nBo4yMOAX6TkrrcyO8sXip0YMOjUgSeblMtSZuAiTwb6TvpTpCqRVwDkFaLboTRlJjRrhWP0HdT
hXKMyaHddSGsadQISXvhHEWWWpxX6Yyf7fBfW7TITJDLRkJlESsp0zxzj/g/KpjMoHSiRjJlGRWm
I6UR9bD3pbC5h08wMJ3A9CZNrDMTApq4K5hU5C3FuXcKHIrt/t9MaYRmhCvjPLVaBj3a2ZZycPD3
EfHON3yv3Ov+6EkIqAZ1wKvXwtCio0xj5VzvrbhCdDixGACvyrtb1nljkyHpWfcYIKZaIvt686Qw
JW9c2m8Unk2/HsBwguHZoXOh+0DhJ4DAyWDVNS6dwrLzTJLxMjD5xBOMjtVN2+OzZvp4+EGXpWtz
1GGBXN7YGjm1SH7NE1H6GOb+20E8U5NC5iWHkoMkEMrZWwI6LW5IFlnLKLfkDRZcc1ONsW55OPls
PcRslqIiUHP1kWv8Eus+Q3STIwmWX2YR/iOLU5soBTo5fomZeJXK9i8v9K5xulH01L5a05Bcq8kj
3ZSwUBYmqpZ7N1Ji1G1hwGUISCMltVNm6SviWjE+7MizawQ2kmabWTEErT7vYGmY6MzT6Snv1jDt
3WfEt1bzsYe4wOnpVpuV0UhRIeZVac/WEL2vB5rLSTJdZTU3LXGeciL7rCzPNZmgjMq9uc2MhTkl
OAI4AfbXbh9XKlUEyU4CsqTO92p3eCb055xKlYooTwAJSi4e5Q4o43f5Vyb/r0dv4Wen+0AAEOEf
clbkbgllhJbBjGX+lqQv5e69fPXZDLtp1Nflhj8V7gYSbQ+6gjqLXhcN7hOvZ2ZRouCiz+C2azMb
4KGP7dRvxc9URxdivBm/fVB4Laezwaxaqs0J7KlA4CW8r34420+RaJ5OVi38PDnnZBezdjUKxPq8
fMrOACHzjqwnW/JO8t2Wzcd2zmzzqyvce9fGwsZI+YbT20n5yjnTxZymWYL+RCgKMjAWN7adbb8u
IulNRA6rk6qw0MACug9zByICH9BfuFPQ8sGaGNykiH06PgRDWLUGX8pv6YjEcBNt9eA4ob1DjFZu
6s4P7R16mGfcyjKM4FN5rCcWEZ7uRPM+qMMAp3Mh2o2aMlmknnpGDr62yWxMupAR1XBkWAiv6x7P
+VIbxUcJ/FFPT0c8y6wUi1Z1eWsIS75uqE7cjxerqtPjGY9XLwc90DTrMMZiXg+lMhjTj96Mfn1d
ZTsvpwCLsAmzPxrLxReSHHnCYTA/faAeNh0/KmObVAOQ2mH7iCTrDtmZkG/WqWb35ngPabAlYs5P
euaIbOIdKqyXi7gaBZgjgeLc1lga+GS5GITgQyiBEgBqAC2L2Yg5m1770IPOm1B3U4DxFR5VFcE/
pizZ4/GroKVGaipII6/p11Y4HEr3soYquAMC34oahkoUeEu69G2pdiCMOfkuTH4/+FQOVSnVyHPq
2ArahuoptsJf0bpOFZgop3bKsYU1uVBoUqEzhr7BWPsp+5Odvv0YBms9iI6Iw7ykMfyNimojkNxn
4AOma2rE1eBqpcq8863qO8AdU/UJ9Vx8arzMoMgvlCJd1imq5z7SZMz+qht3AHGia3tMpvfQtPqY
fwjOrSym83/KrFfcgFHMpKehyfR1Tq6QLA2DLtb1Lhnze0WHcb4t4OAHNHKtNLWht8sQyRGanZ8/
SNKk53x4uy/XS61xKD9JWp9IGfB5VepZl9eUAlgPegTbw4anSz64h5dQHyczfN4TLe6WjwkOXJm8
1WCQl25JS/Oqg2RsVqZ3i+H2NbXpI/loAvttgXznK7c6ltFQltkvLqA/9EBuze05YYCIn9dp/7EA
k6tF6ZCjzGBfTeBdiQX37qftkHs5PF0/QJRnW4FAs1DtEmYWC1x0/v29lKQsdzpUuRSpdogv6MCD
bZWdFx7hlNZjCWziyDTNlH0D3C/D6dPpYZeVEkkSlEW68s4oYUN/p6UWNqhmFKo2vJVtyYoR5ntP
FDXA83Vd5DisC80kk1TgjIlh/K+iHqPcYIp9s/vWbOQWLCZMZyQcCuwzXTmcVofKykMzWArnYSoy
FKL5NuK3x+UL0WK3C2pTMTsjoGbIxgCbQlZY/45k+jgQw9oDof6NiMEiJlv0td1F87jSa4T8mUaC
oGpdvD0Gds6yG8sMJMvuEvLtfu8HKVmCv1VdMgOUVnxXaHrz23G1Y4Q3KmN0Cn/t4Etajav2G1s6
aPvc2Us/eWVoQLTZ+nLHWoEsgXBipKA4IEdEGe4gTzOYrKSN2rvXt3+GzMx0tQxr3J/rmfF/JTIm
2MtNyOR11a/4XyCwBpMaTmxHfDhjf923v1faHcur3tytjc8bKb9Zys9Za312gXEEzei0j6cf7TbE
SPJGE6Ax/YzxVC9Gj2FN2bffNqkSe/sLFQrXLCXJP2yQ7TbvF6PGTH2ueZAcPd+YnWSjtRijjBfg
J7PYszSyYjBSSvS4RiVvWMqsPlrLFIswoPNsIPElTvF+B/PUNGJGb5/aTur4UTcxgqyugiaiYsWZ
UsmeR8DijO3q3VMaYEAfvf1DGJv+4BcwAzc5UahUJPQiWuuQPLWEQoZXzxJyybvt8Nc/XL+E+H8v
atozGoczc6+coyoTraX3cXF9BDUl795MsopMdzmWvyVpuQVt/1lkn4qS3jYQ0ct6zznFuSUBBr04
evLKvxQVhIzr6MqvcUGYLJzPhtBs7oHsAoteW+bCpYFVgAbWjKxf6/6FUbGZEcebDaQtvsz/fTii
Rjbc/qrO4Eavhr6T5B+ECGRL8B8olI2M+O8LkGSgm09K1NPJjXXwwNh1pab412iIMWZ7L3C2U8ns
71qY1JDC3GmKt3RmKzOsJp1rPLUpIG/CLKuIvFIcDjjtenHn2w9PFTIYhgUn46gxuYFxS+BjRcJZ
RHWQ/ZW4sB59Ose7rfjONTgL3ILh9kMdmrqTDdtJ9u7DHG7tBPM2T0PwDJuG9LwceMM809ktY/VZ
KxehHCfiS2T9duxm/i4be299T5wFAVLOn9/Hkv4Naa/O+a/k64TDJW2qqSbDyfA2VcRlEjOooJVk
W9DlkBjlRoenTd54TGU+HGo+5glJ65y3qrQK4p6TkTPjiPkGmX32103QKbsNssLTTHRAMsco+qxJ
q5AvdebA45/cs+6i1igZpfv5H8s2uDRF3zO7NrK8nnugPjvbUeSWNUeS2wraoPhAxXxXA2Xxj0CV
ncFKw9r0YhFlxQJD7r8K8o3zxVfVuRrsiZeTGpBQA25G2c6HJUZB63cjXKB/ct//Cq8N5WC2ww2n
LlDiju/M5ICI/fXu24Gao3aiDUyrc/WhW6eyMb8hOqKWXmsYCnVdk3b3t/9eJEyn8jS5RvLvzY8u
pWMSk5X8SAvrlILS4fB0kFsJxEyHAr65/XPsOTOKKx3ofIDF+KOou2OOYAAXgirrsAGERwSFgg/F
G1p3uSYrWStRj0yKZ3lVegxjl5x9GER/0WZ+IR6/+/aGaTdDqO7dixe5OSBpnfTdWJBHgE0YiPE0
A5x+nv5UTIEo9bUlUR04Gn236etE4epnbbVqOJGAW2H6/MPA1LXQyxAQHtNCOUqcfW+riEbDQumB
gueXd/X8Rwv6UdSAv+fA17nPtySlWeuNCnmLlu4st3kvPBtOMNliSYAMyIShJPG1Y8r0M5EJjTDt
pdudjoWWJg8GenrM30ny1O5PLleRDZOvBvGaKBD1a2bRVnADt/fEktxzwNEuIisaKTX22bc1pL0S
Z62pVrXBQo00hnMrxyf0F5dXG/TWUyGNz1XaO+3HGOC66V2DjtVfdeOUiXSUDY/HpaY3zjohyh6+
z+OkFLNBZtE1wNhufLliaCQ4Qr/4Bge1JjILXkh5FhsaVz6NHeBUrHdpILqV9qnoJ8WZuXWeEVQE
tQpiK4/SqUs+k+kCPmzFWj/mX/9+oI9DZVborzLVM1/o/2yGxrwOymBWfbjYs8Ju+hfPw7+BDxeS
Ow3I67em3fZ7uVrftgn/UiGivTcVcwpPhocUniQQuxHYpiHdv/xKks/BVLEWYVfTSYRmJyOoHsN4
JCu5toK3d1boJHr4QkoFacsLFa6PZ2QdOxGeqC5crJXpV19EfYOQziRmVMKv2/easQ7IzeI2Ns+Q
qlhzRJ1fzzl3tqstKXTRxPF1wwlvFUPb2mHRIpm9XllcYmFvXzHrRa13fCl8ygS14pky+Z4vbsSm
MXIZKByqUDXfRaKqrNFJGh9RW1Qf9Tmin2PnYly470D3M+kacbBiKz/29iW43kcIBToYXcpinEYX
R6DrhBV9auKFFemtsm2jB8++v6BQMBBnDlT6ZcpLTExMu6aiRL9sqxkuAUQjIpVzUUUgSfo9t3vw
BeDWdyjit2m2WIxlsFVGsUYPGAddbNjHq08k1kgzwxd21l8L9B6iSQoAG7nliOCUDOo1+0/im8+0
N5fIeENy/Fw/Ky+iQELp7+bH4JKnBxH4noN0UeSXBms2ms+eXEl7qvkWTfnbzVgYo680iF9iLXhX
WsDN9g/FHtO3y014xN1Ffm4wC2gWjv5Uyr0s8ricBAJn6fRum+WyGn2U/lYgqkVNSNClX/uB1F35
TymzXzuH34zNbsZsLrRI7GWfAlgAioOkPC3gdfoS4cOUL6d5LswCo8ZcdK13B/+C6VjM50mkwn9f
g2+ad511k9pqq7biY2CBWGZ01OPCfveva5ynEEVBPJqzsWENimajhYxco4Powlsj8YbnXtzNJKCG
QQWrD2tcxFsCFeetVXr9OY+FYW5lED63aqKIYhGYicCynzHZh0mx3rp9yKthLeMZmTbah7D7dG2M
XSw62U7ozlMALS01ZH0l80dwdiOWBTFQjWyKsJT++4mMF3NyW9Kq3uiai0bsJ2nCVySo4Gg8LECz
qj3Ub1RCsorUIRq9iRByAxj3GbtCEEg/U0Yz/9oXVT5Gj4iGFiK/ejWh1RE8FVUiUE7QyMp+IrSr
Sj2PoTZLE4CX8Dx97TQ07ZG7mldd9PS7Pnbff2JSM1NEuU3qbVCX1cfylfGC9g1M6Ooab6Z+Iw1Y
MmsUsjW+7e7uCCcgQ482gqZXYDLrYawFxBJY9lgKQ56WJxBDBDnBBhr09Cnji78R9FJEfL2ADPEQ
iT3SpPlWG0O5qCWitiyKSDLw1fERxlfJ9MFFuWvZO8vewk3RsHpbJO74TcRodAdmiugP7usEgATx
pvOFMniE2xGHoq3wao2anmgd3Aug6l+BiwAa81Fwb9bSlvRDybFMEaESEEH7kSY8jtZX15XRpo5a
qLhgJ41vyU2Vu+ff8/nFfeha7ScO8TSqmUYkO6KdYPQnqOE3bh4thPfK0JFU7kjMwQmXF0mBM6E6
S0x0opD7trKt+8Ja8LoYf3hCS1ECxG6UcvfOvq0wmX3sA6YYa2DZLLoU1xqJPdaQMJ3K74kJdkdH
LQRFuZllVn0P1w/AA3EZS4b4GLsFJdXYAo4RBNcAfbINevmvXgQTe+uwID+hFeGU6XIe4HFPuaUR
YaZb8kqqPp58UUVd44vrUC3lUmrFUrkLKWTqhkoq38fsCndtm5iwHOBm1OgP/xSo/biwmiGZaD1z
wWEMz7iQ/+piFDnROphW34JMvpmU3s+sTkY+mZVPwwReu4EyPWqEjeecwkMObgIWiCGQ8b4Y7JoD
5U7Junzdn+jsOIaw2rg2ST6Jyd3cDsVLVgCM/vPEZa5IPr+KLfvAwYefqvEPuClkJK4x4L4quUmm
LgXIhrbuwqQpjKpZK/a+APTIDsAJ7nG0+UunZ1laYH7p1nh/raxmmf+nH/YT0k+LZztmXt1S/xo6
4P1BU32BmKT27046nNpVQv+KV91gcPKEEri87Y5p8XLHRiKfWAJPnP7DG0V5OF7+toykAHzai1n7
q5gqD3Ya2yHype5FvReuESlbagKkK6CI7pqrKFH9mpIohbKklWpteQnXMm3ULbaju+eMtul+pWi4
5p0YAbJLU6h0t8wORZc7X+PzK7KWCBV60O6bjvYFvQ392Y89fHludRsSn58A0n9vyL1giTizUpke
dywm6htYd5CnWR1HupI8o4Y39mfuxjyATIoxdYmCp0mQjgBK4K5q8xThPp5fV74EFVyDuQi/IqCe
LzNeJwt7uQNDvrDfYPkGtY+asP/2Uo/v4NFTk3XCnC8sCml1nNl44K/+yUE2Cf0UgrU60os/9rd8
uh5RoXah9lQ5370+4HVkm8fjA2rPeWgvmwn/4AMBtA7ss5LI8CUo+kgLImcvJcnx9O24nFIR5evz
WtNZscCjH8gcL7ChyeXSIMweU2Qwsd1DUtwe5d+dwrZ/YsCtALhWEljFYsxv173Uu/qZPK/eI3uB
0TnN66CjbGNT79lyXrDpHAVfDE1RlAWMl9bDzrroHD7gnb7WzAa0wTEC1oZMLXZ+9Z1g9AZqeZVo
GRLiEwdgyBKGMnmcoZoIPE8EEExy8If3w94miflCyd8nf9F3iBVnqS3mS4SVI42XlbtrrKgk+8OH
Tijc110bX7MRDnmMDuRUBobQMHJz8d41pistnFBCxrtZPs8nqBPNInqKYBARqWtZGMQIdukuvoA7
eF6YrztZ+cGebp55O/SIaEZs3KjbNzURyDRWN5EVeH2TJSrtNqYvSbFgDrutYf8JDmyK4Ceq2irI
4E7HS1wDBOMyGRRkFEYic0qQMkwnLJdoPdqB1QrEnyaZ8wnvwRKM1qpLkMPO7OKNja6aY7dvk7MK
CSi537EdDs6rIX21VuIRSBb8Gxh2GhejI0qxIYtgl/a9CQ78k4joiePZet0V1ONXrlKMV5frLd/s
1O8oH0j0If83oLmiFLzJCCmsFX2z7BHg87LPJ90rI96P9UvmuvAXTvxeey/t2sYVgu87N/sRacBw
GyJTtBRMhN0y9DDzzEz7lpnhD/SidceMuzqfRviFoqnRpqAbxS6Ah6HA4vIToz2mU5H3mWfvJFSi
w/d7efYXBJqCm7XRJXH1DLG+MLLdNVC9ZZmREkp7NogOQGNE1FM9ncuj8aMJe36Pp33TBgS+wxgq
ATiBbzidXbupkVdN8MIv5ZdqdCC6xX8DLFja98eUovkjrreMg9S6LxBYn29Uku5DPrELr8BjPj31
4EqWVu3D5KNND/u5lTHU9C5Sv2QqZnOhz9qkzc8Q7NGD/g59NKUFux3pdpZF+UyoLeR8td8ByYq7
h2JTM2C7Vj1Ih2TSy7+a7Ew1bmPgqJujuS15aQFKk2znpceGUbROnRCwxsld9tjb7fEAUGlYIvle
GcOkWREW6RQyAkq2dbQeL5ywWu1FsaByPsQzJhjASy9HoO6j794FiKiHn11kaeCPr2ChR0RFwJtD
OwcuO3klx9AAmWN/gQPy6SfJODBOyyEtBnD0O7GS66I18plc4GApRJ71xkDuWbHjYJZFRz6sqq0U
PpOxDaOx3QfpGiShAvhlyT7NCON2AmMGHUcYDxw2d5+vrlqpQREiHPukAsCOzRBgBk9P9zIbiJp8
+e29zBeGj+6vppyCQzQrFBka83j7ynyKGNdc81mtmDeh1vYGFsmuyhugdH6HCM9Z8Fc48SoF4D76
Ox0OspDeZJlzGfOS8HtD66ZczZdN42EEEBppTvZiFp3qsHw91JYrVPz2obJ7X/4TJGYAidhwEBc2
LvRn39jBHQpiaKLB5OCaLtZUZe63q9yGaHAIU5E8RuVSY8q+nevqg1LmFMC8WMby0voOrlUz4x9X
DaGfX1Z4Mf1BJBlWSKKwpXzaBMnRdLvMiduuH59CxlW+aWLFPZA4/oQqm6iviELOlYsPq+9CKulk
iTfkyq0Z6ly9P+RF8NRaS+7il3PHbSGzapNw4qpKn55Sh/vTFl18FBeTJ5oj2VYR6IP1RqGBaXRS
Gs6AcGlO/YvWPsVdhJ/OVFuPRrh6+cucE7QVoM7GIUDi2LuyaHknp4/QvqBQ76KSiwAtmEzKVx7I
IoE9msyWqNMx+BUnQ23l/Ktv7b0d0z2rTjoWIoOoIegjZNsD4G2Dqv5k8THSzxVeNiFtgYmtoMDO
DJvVKdY7OGaAGJRfjEqv2BKfhrMnrw43dfv1Ys1UBTCJWwHBEPstS41Cfd7tx1sXH8x8isQaNQdN
X8X5N2iYIwLtnx2WzX/Qk5rZ/kn/f7hrAtlHUd2N76EZlNq2HRT4FnuL8xaNenhmv7hdEg/ROe83
9vTda9D6Az/+7ieWFVkYgFzYIex9DQv9i4KInIB2WRgv68+CW9CdoLUa2Y3U9msVJ1TuK8YjEkK8
R1QKAELfyL0a5Qc836+glr1IWpXMks4u3I0XKIbnPhOMnspOujgroLPCXZCNrEU2gqTW+1VWVCrG
70GcPnmxDq463+/KyY4BVYaEhO6tx55gE4I6018pLxIVOiCbD42MSn7QDILvmJe3zcL1PiIHmIdk
17NrtFyA3AG+bqDGO+0Q4Z+/ISNEgL8TyoE/q7wYg7aVhYqq5/NFUFal28aJsgkXa10Ql/Judask
fn3oNJRmbdkpnLWN417yfHkPUNraGtSsYv5QpLLUDHLrOk6eJ73yWQa2v6mOREz6xg89o5UWjbRf
g2WOboo6HeT4e/7O3W3pdlOq7S5ETJ+4u8ZN2BIrnbqJ2X2nV7NMM0DiWEmlz1dTIhR6WL+IxPeZ
nAcugEL7o4/KXk62oPkf00ixTaizQ/l6/CBjtBizhVzGq1ZBWRmoBK7WJP8Fb47ESR9WezuKC92v
agkWD5pwOJ8L5P0o4YM4FIA1dR+eopRAMnwFOzq9Z6MJxI2lLV7uVjyGHDAgp8QQh1+EDgyLWcdj
UhRdHFAueZDAG6dfbFfI4W5OzI2nFKEgcfYePa70GduFBf6CSjD7i+wd6xaPA0YhumtXjg4l1zwu
KvIe04dWoG/OgBayqx8kD9fiXpQasjnkz/WLb5cMSwx7rMuq6tJT6NWW8CdPyiTU8jYUwWfsENZO
XQSHRqxJeH6PJRVpXPzzCyHwFLVew9QIK9LIqio5B0c1EE5TCcYJkYRWk3yevHsa2ZJXonCbvKm+
9MK9voPoGz9oDlQdW3JtoquJ9LEW34+uJ/+jgWlsuhI4lBEGEKt++vZ8S6x6aT2gEIpkCGBFv4TI
xxuObpJJ4WgiEdKB/G2yAuFy1Khuq4JKYFGfu2YhfjCh+7sjSkrhLbhRCp89NqDKqx3jvGhyrcJU
FMFV2jVv4LfG7huNYDTQR/3mw41B22fnWSmn6MB9yo6sNXUbBJiLU2DmhslsqxMe8mB4lz4aHtrf
XST4/dmyu5gQVeSRDEdJjPhPrHvvkkF44EPxxVJbi2fzaf1w7B7LRQ4levgXrm4ThjO75+sCvdDG
mhgBRm7DngnNh2fj0Vn9LKcizOueGodhbHbhndVupkBEAqGs/ajr1Tk3/r19g1/Zt53xfJwXCWtW
qnyk32nijhzej55DvIkLsP2HnSyaPRzsURew0ZdvAUW8qyo9SlBxV4jz0S4XLSjyPXSHDzV0VufY
vNvAqZXSGBqEAOmAC3x0cOp0ehw/d97UUHTKmFFaanX54OAs1ZrQE+UczP9HGCeSr4cDRoe663y5
8OtSC6O54NwKnFpAtFHcbBWzH6NjeamiArr1GlNJHW26AUpotSCx3mx8IXPd1JGvTTy66Piz4WjA
es+X+ti2M50Q2BFstISNevasRFqDSOZzU5TdBbXJSwtC88BM7zQpXQDtYG83wQiJd3J8X5IcnnA7
a/ITRUH8hZB/xnC/jUcN4rtdnjjLKehkkDbbcY4pN76lqk5QUUtxXHWaZ/fgJC4J9PbEvfsaay9k
Xj2a+WgedoV3cs/W6uu47YcvoWd8qFCfhdbjNBMqfLbLbsJqGX21tKn6kMXw4xfzgEEdl/cM3DF8
tuQN9x/VTSOe15cLSC4popOGcMr3pyLvjJd9mQknenJciyRU/Qki+geFsYfrJlV35KFJ0M5sR/0d
kviVSJMpN9kOIAWbicEfslMChU/7VgkzzHXf98zFmkPseANhbdsBl+XIVrw8F4rOMni2R1aN1u8m
iMNjbq4J16QOsGU4gzdn5K7G5EIM+7+Qj4YD3XsTsQ6EEoIl10/tbWTyHZiWoeyplMwrmLt0PJQu
gT32we2SsZwrTNjzw37boufllLjW0hwYMOmk2fFZnxbkB/wHi+YJaKPueIxMfn5BSiOlkwHdBjt7
8VuHqkCr05yz5RC2QldwXmFLWyN0zmvCA7jTVDX/qkgq4sNvXItQ8xACJyJpogLhBer8aXqX1qjm
5tNUtBRWsBeO6WOR2X5gcBNLXDUl62xs4EPShI+QRG3Omg0TISf7ZVz8NMqG4xIU5MKMhSRLZc+E
DGiAes/wLKbAgNvVy/2bpUE/HnjPBvmLBHo2hc5yoF09fE6s2ed+6GyMAgKA3zc0UXpAfQWZrwN/
ryjmwtxWvMaNi4G6o4ur/fHMLkmua0HbN0n+jzKU/LYBx0xXxME9h7Us8qdIVLGx4pQaX1Xmuc0w
vYDjnR1zXq+uYYCqDhckzJdVhgRxWTSyOwlTeClF4XXVkhidgpVbLHci3F69CqjqP5H5TT+eo2uC
4dAqsgHoK8DkTH2Q8FVc2pCjgPqP/kTjY9lZVdNwMnNXjrfN1Obeotgd4KlHl3ymQJQ+W41cRIN6
oL41X16a/C7sYAAvYcbSGdIxZrvm1Wld4/8VgoU+EJTfCcUZeqNt2qyw7sBxZJWkjRkrBnBEKl09
Z87Slkezmu3moVQacTXA51QoKHCox0y84qyD0By/RnthLYpD/HM/5Q8TgTKvEB3WLgi0KI5SQvpD
gN5+oPC+C6BpVcwSz0xE5MjQKCJ0gNdNEfksMdU3TISn+nTgUdBjXgXQRQVEd8HBgJ4mVPj9JQoE
Pzq3Tu9MAywgKyuetuNhvjulTRlk1KSI3a7yaRizAMp0FzVeyn2O/d2Mu6SSTR98/Pan5l1x7J7G
m29Ih8lIIS9TBq0J36uabSjgMM//utzwzUBeMc34pQi5JF5tRV3W1HqbeR7ZEs/+J6qnSD5fRucI
F4rbv73OWWZDqnmX1fPgwlGPDG2o34WCQUXUWI/EFlAaUZE3Pj4RM+E+K0Tyy+t0EY0SMKYHgnYl
kMDciFsYmtOfFWa1CLuI11xpC28niLETa45WZn5sHmYDQ4YS+QoKv/yHrXT/PScXCz9MHNJ2Vgzl
DHCWlSPr8B1xQDoJTRBvmSrEa4+JP83uR2huC3STTOZqCn6eNJhNL6pGg6Fuafdd/XbloEd5nIT0
fhM39/H9Q1xc0g3AbnmHDIlWOKZSPwFHVxqdSL61w9eJLeaXUOaFXvcu0G9yLT4MCDGcsbj5Yxpg
uxeToRlarGsZPztfmxbPosX7c4v8Vlw6v/2hzIDKtH0XMpT4RnBPHvdKaJnF6H1bltOEdnLAgRwz
mD4j/iGoP3U0+c0Pm8OQKUZ5Ft1Hx+VctuPP81LJ9axdF7H9l+L03aDQUux42o9DcOYaSAQGTfm+
3h5bn/FdWpqhJjtJw1Zr5rJBax74hZLseuZ7UN3ZQVSAZKO6kYMeYuanbxR5Me7mbVysHqOsPB8u
mptsxqjo6LjebkG211ickQf/KeANH9cZDPVL1va8u1jY3HNhyM3r8lc7nQ0tONZNN+/aE5hgpKrX
KXZlAkdzJhesEVaSmybkIatqOJSKVG21+xv6l34w+jWtxw/pP3RyxZZEis8+458U249XAx4FQ7Md
HpsQ9WgfLOdMc4QRb1IdxmUQvQox3FKgPKOZXP9E2T+Wmjs5J+g1Aj3K24lndd+kxXlOh8DwNL0o
0+ZhdoyOgd2RCeuocaipZL4HjYb2Q3ykkabzp6v+ogeeNzQXXTnYaDtwX9rVUeVorZOWbCwbgtgN
9htxTjHs8k30kF58aTijpe7AwC+kezf9GjnyaZqdgGoahuUNMm0eKFycLLp38YvqMqeUIrA3Z+aA
UzdIKoMzbSy18GpbzyM8WE6ib6Z+9+aPdqs451IK4Z3kQpUE2A8wt/TuV+qNJqlLFjj2mi11iI3L
dPzn6JUuXyaNd/u1BJfEQeQN8M5jSxj41lum++ufUJ/t6/EjSKyqbsoz3XxMq9Jzb7Z7znBVjaHY
nh9SGl9T1W8YTy2dTD29mA5qldxyUchRljN3EfeH5pBhpQT2opKPu+5ntM15JGjXS6gsNP3gPZp1
LrJR21CfUX70SjICs2YGbWXzotEFrpxnCRmh9GFnwKibW3W4eX3OnV5YWfnf0vgqowM09QH2u+i6
v2MjyBkyRuxWm5g9DfAQpe8ZUrjedEmblk4Rsg7o2wAlvlhjAcuU05Pj77U6Z1h6yo7oaCmsYe46
Hyl8tp4T30o54PN3l2efJGHAKVG2vUNRMAYVh03FRj5/CaShtlvMVaDm/7oyzbaUQJfO4SOzHm15
+w+dEeOTvtihxXsqf1yQ2El3CFtFkGW425DZ46b+zjmtnHANECQbMrDy7Q4SlpCqioJITd209rM3
fYFWzbSUFXvXNtsZO+onXjbHhnu4HcbFC6VCe5r0ZJsCaRE/KiqB3DBtisZ7agk7e3tNFxroV1UQ
PRPXRiQj4lp5THxet+VoomgcsmppPIcmtlpeDZe1DNIvsSivv9OEb9ofEZ+ry8kFaV9kuMrGG7XJ
xVbWKsQatptgLoz8R2eN921+ZDnF3lN9OErm+pXKM/uUlIwxlF4HxOYmbHGbJ7N/QPO1LaWNa6w/
QlYZeMK0FuFESIGT8YuCR6BKRuBGvnDWa6jLanmY/rvaeyGniAsnvNUXwurvxJS4fMAHsfncaev/
ETpHEol595Kb7WUXXJHAapz4j8RF/WRMqcBDTbcZPHlfL+EkxnSeTZXSbS8GLr3uic6AvwBmo6r7
YBjAv3NTQo+Tk51ucxFcacfIWm8cRZANr4POVvvSG8an1yaxQXj7iP/VhUTOxS1HFHLrlSTbpM1U
052bfWvNcKpvCqKVILLjEmcEyqVzxzD9poiqYQHr6lCOKjmME1vo4fXiaGs1V11lrSJ1kMOO+z6c
ncwGuSDozXgOmG6wggWC54qGvwoV46vHqPY9G6SuyNOhL72OK2nyNtVfDtwCNAPm4ZlNBlj+NTNP
S8pnMVQzU0UsnagQkqkdIL49fMpzeNkvhf2XeWR3V2s2n4ovtmUnGxijzbTAWAH/JpMls8wcNtW4
XjcIWmvCDYcpOthFagwgpY+VcONp62daNqYk94GnSs3cYEodw7r+tV5P7xHtdN1WCDd7pCeYi4fZ
sIGmdls70+VRRmuowM5Eg1Xplm8neCSpqECujDjFiqTHMUHrgfKNEud85A/bLlsSU8udIIPXCDYm
R9Ig02bZm1gpRpD4vjJHzhjoTclkvaRzPC3O96C6ZAFt2lnofs7vkJchPyAAt6+TSaNkqui6HxxM
H84jtTXHgm5lx2A5iWmJNzrLl7lzf3Hr+pKSTuMaA6x2LemfwXVrqtRad/Qb5J8pDPT67A9eVjKN
3ZCFxcFn9gkoHuzfYzrUF2lnvtnx2laGa1u25MSjYfER3WPnnFiEHtkEIwEqz5laA+t9eWnApTZo
+UP8ltexbOOVlJCnTlrh7wxYzJE2kfWqBXR4coBZe9i4t7/Kv6ZlaTzpsH3xWBxUyWEbYZE955+g
kJmzPv283QaGxYkUvEuR3Oi/JOYAG97bfsH1/bnNweX1D3ZWkbsKtYYuzcd5HuVL0oU5/p9fL4Q9
9W+pkHUT3/etD49PBE5n0Ie91C9YwncPeyjzM3x3OrdTKad0Yucmr5bAIKXCahtBRdmlsFXe3Ntm
zESsb08nT6TIl5FmjCCKx9zohtt7I1LWcQXZ81NtfOzJ1MzxN1FsaEX3gCoBimFcJM1NMuCBBmiE
UC4mx+aibr/2bdU7eyUBu51jv8ckcXe+TPcwbvvzVo/Xf9WEMzA5PTHnCS1SynNMHGIt2A/gxgf8
xhO13kg8YiGAEt+BDYmMVRYLHtc4yC/3Bmj3VO3x+YssQE6+XWuMTwftU8lxkZ4rsFCWv4iq/v3E
sqPvfhrj+QqlHj3RQYXpatnf8LH8GvGCiNBiDDdSXUUZJNPACDZCHSqIjKZLf0aCFja5Lfna+BGZ
mox3gZCXbYFgbKjqtE0XnJiQyH7gNPR4u4fWxJDmD7MARFV+/vi4JGxINxKVqr5GHgeDTv2yBHLQ
+tx+mPedwO07DYtXtKpLuUeaQ54RHNUz0wLfRzfwPw6FyNMTXOxEzEG1Mg5WqsMv0drpvU6OW+vf
LWGm7mdJC7Ch95EmOw0wC5QmoZjc34QXcjWtM5XCeFwwZlJ0bxj//IR+8KtYqCCiSKnA5hgyl1LY
rPpW/M0ZNR7Y8lW00QQO6WUOffnpa12xz+S8kQw+kh1fFuwKsC6Gv/z9qgWahswhwIQ5+TPYKZqB
OeVHZRC/u08R4atSo5T1ewJYbKWG4vF5XqOrdKeDM8MnWrl4eJ6rquQ/fQFSttg2/uzFzBsmN4KZ
AF2/VaQEn1ALTyqb9F7/U1rvbicn+vLZNuqoOw7W5kYo+xec2sjGqODz4JxFRE+eEqxXJUsz2LD3
H8gPAQR1nM9SsKwvqWzCeqYPaSFyIxrvtaElMU4ZypB18rzmQ2N5UKu4XqoFGw9FAc2NUHD2bKzo
QGnI5xqc7wpSOAjuBMbISQbN6ZV7lQ9lw2UpV15PzdnFlpwYbH2BJKh+3E+2+JV1taQ++2S7fgci
XO8JsrXjOGMIblTTzXX1/yELCDxqFNTCgDmFQ2Bw/1CuTMJNhNHiphwuWHApadZnRcsG8EyjugpN
r1fp4WwWCY/Ti/3x1+tL/Uc6nBvouwG46qFFdCe8WY3K9HFxp2r3gQ5Xg6ANYdQFl+wEEl42V/mH
Wk6uljFWHO9oatzIP/jseGm5lVPmbf+Ef7X2GW6GXoxirQyqi5tYS86Pfpwkt+nb+yTMMjfRfZUb
yXtEQH8JX0Gr+ommpux2N8bwAJ9uxCBRZYeqrYZvdv00myOqJvEwezxrNXkdBc3iH4m8k4kbjOpj
2Onn9AQWqTiq9W8yjCAXKVKeaKgpqr3GkIeA/baIS3qhFH27mvapeqxXsf9HpnfKFtM/YXIPlIkD
Rw/kYQPDdLFkuie5fL/kLLEExDr9tL02Yh9nBJkM8WJT2lannGeGbMTK4utAZuhwmc2lwjoEajuj
jS4ogPUWeTwTT/mNTmMD30G9hFXcAILi//9HRWCD4EttZZ1rO2vYQdgGaDUmreZ6RNww9vwREwM6
HpaUOYXZGrSOieZC94OC9j/QG40D/d7gcDfvAEYjozgOY8m+Wi7LAvMyIQJSq50c4LuI0zQCfgHj
+wrt09d+x0dP2Jcj1jVT3mVMD+TrT08RwB2a2q3FY91iKt0OmwiF4431VwF6IzE/WuaZLAeIMVen
yBmbuktu4nzVBjp410JApBbtG17bGSqPUZlv+k9IkbjJuJVX0MrqyRwj5D8AU+2leC6j17O7tOMk
ZCuxjeANseXKPOmntDbKfK6VGNoTLJr0Ix7Yy/AHLial/BvPBVbORfW8RNyx6k/yJ9tH9ddrRbHW
z7fNa2ZKQmBnUin7JYXeT/Y3cgGa3BIvC/IrQEm6U/gBAdVZLJ7aJ7LxWkfglmi8QA2O/kdLwL2t
jWBPcdg4hhDj5xiplmaL6u5jdEAtg+JiWNxHTT9T5R0k3lCJha8QTuO4um7aejDLrooIkb0ml8bv
HZ/gCXqinLqwCosyXcFOH89es3QLrMHXdYLUJYjgwDax1+4CuYhQWc/ZiIcbLCeyWtBizLZw2EL2
YJQ9k8l7HD8cM/x82GAuyxEJ4dqUtcQpyrwmEs4MUD7rUk0kDLUJPvkAdPJBVjfKzwQx+k+kimlp
YL/6BiSp30cBhWcMNpM/457/CRecnVYDn2ZdBLbbxgQkB9rb4MFjpGjpOWX66JE2/td7tdV+RFul
mc/3mNRmXQm8903oZXDXV/GpFcq5+364SHC1eqGYGzRXwthkZWzErL14QmdJtYBD1RuDQRdkYX2V
Bn1uiB8K/IRiondq6+ossUIfpJYVaSYKnaAButw2+76Ey50dNCOn0u7VFePG+2C5ZrDGadyHf3bZ
xA0g0L2qNSQcE3dhf3enY4jl2qNDS75KzcppuaxQIlN33Wk6dbSajB1NGz92BSEc2qaD4e3LBZoY
24RikD/8x44ds2Eid0NBrEc+squ9JpkiFOOrvKRwoehIcEWoCCFJE+NaArfVjtAssMq6BapvW9f1
EeF4B+goJ0YHZcIuu7mE/ONBLNa74lgLVYW85oI4/6KBS0ZcWUW6YL4LGdMi4WbGt+aPrVMkDKJO
HDH0fVByH/STKfMAHYV696lMw9H11jSSPtGSMOuNKZLZ/QoGTiSK9pW0etxBQ+VcPVQNXG7Box/y
s1P576MhdYRbe/fkw3lUOUbNatjDT1TtahUS0zBdLa1e0nqkEErIy+MKdn37Y5DIbB3koOkvKsvi
2PUYkz9OPxwxy3e5Q84/u2xN9PLmFe6ivUSpHfmohfhuw9Eg5JHHDTlvL63ZjI5/WKgzAZdec/a+
mw58J4ZkJUbb3yT0aHfHlqZh0V72St7f/zp33NC1iTgW0JWgj1b0tO23i9c1OjxUB+x5WMGFWPBT
HnZdsahNYQveP5DDEBOOoIoXA5DNgJJu36gD4w8mdvCW6NQvwvVDaN3ZYNnMDpKZtpOaN1SENbwl
FS4XsUGVi9UCbHF82xnDtiwNuh05va5eFneMB/GB3PoGQPl+mYrt+lIK9H1AQg9Qw95U+38RjgCR
6PjljfOuFFqVOXpgMexRVc2fhhOGUAd0VMlh5QdarzpHf90JobYj19OZba+//dPgFqzl5YrKrNDA
7azFyFQ/i/U3jGQl5ahifiwWHSUAhbI4yqA/uR8cUOitabs2XsbyflwNtPx6P11OF0KEhKlrqi5b
74DVNn+Sd0+jeKJUQGSfpLjqU66nLN9xkZIFlZF33prMv7szvOI91b7u3zTep4Aa0o23y5DKfZ4c
K43+ZqlZ435kLL0J+QWZnaU+CWD6grWa7w6fNR3POlikgTI0ZWxyzQXbptv4flz7FzW155pn24EK
zhilF/hX3jL6+cMgaWYBfStbyaljiu6krCfp05r38/l5X0i8Yl+o1+5XZqvAB6t7+mfdtEgbv1Kk
eHKkuJZUWNwJ3D6jO8sPZDkAenvOFJHHXeiAY+L7Rb1oP90jzrN6Ireuekek5zsODoBijiHFJD3H
gn0xrCQAMW0wwx/mz0Cl9qJJ1RNQBn4mt9J8VLFRbW/aMc9+TDpLTCveKOMxfmiWH4ziiU1DMvgu
jWY6cNuedk4G2m71eELNz/gl2v1u1fgFv/0W034R9XEWWwL617wZJdMQhdw15VWOhBg0g9M/aPI/
hqT5E/ZTiIlolwsvT7AbDj1cNhRD5jrh8mwfzYGVpV2W6uP4jwrSw254lh2QnsVACCJj18/1feP+
EWcWXbx7J9qrUX2X/1OJt4K3EiojDPoj090mcJ2iTbIDGJO8TdAtbjZrJ2SV6Ncn9+U52myiZcxb
tvmLTkXYeh0zP4v/25V0PPOmIqvLvgU8NyBvEF0gEBHaYglwWDo9PbmH/vnw1oR/BfNfaZqe+UeL
knbAAyAY14PaqcJzmT53bmZCojzVUBEodFjeipdezIM2+I1kjpsIGIMS6jBLPE7e8cG+5XCQoHH6
qpg5Qku6TzSWq5kf4KS2yJEPMvGDfdmnforILGDwmUTOpDXlMrZIAokJNwZR64jbIcDhyYtxdVtG
HNPrMRkvxLI+Hs/GCmPXyVmYTUwNok93W9+F2BiKieeCNvndfQyGL7//YZOZfwENPoEBrJdLvKWG
TbN0EaLVOEOqOki/xUJVkKlywqGixaLToeaOdgS6DYxvxyGQIgiNMc+k/FDvgBJ8avRb9JDLftqx
Kf3Fq943t0Ie3+WtCwXp2qJykOuxc9exS9X5bU3azcYYWLVNNtOJxeWzQiNt+TH4z0KxgW0Gvs20
znytEhT/FRCoyJuORg1t00Abo+KilBLV3IrOhH4fWyBUtJrKh/ScdJZJ0HRyJPlLM5b3JQO7to9Q
oVYV5qmZ16gMHx9dTO22h7XpKGwgUTVelWlBfWNn+ivajEMtttW9+ynNj94sd49qkUjYisFiJ93H
Yvyxg5n19Vn0btvZcRsZ6E2dQuwDQ4dWvgFsaO+nvcOa1PlPHze9Hlyfq0mTtcup1V51LAmtGGms
gFw+mR+YAQfgZPaWej3oyVDVRtnhE+O6y/z/bq0OTbeiuctYuGMqN3ta0RKOmLJfbkxzj4TbGbLC
yHJNWF0z+FRpd6g+Bo+e5cmV88nKHMnBHEFXDF3goUxXmqvH9KysuugFMS3znQgOuWF2WuhhPyZX
d3CWufxXBfrFPwAdJbYK8R2QrIYT7RLm5qteu1xtAgaX4ZZh6Nb7rWCHYpFbssvJqkAziPUyFcy6
vF6q2XX+MF9pSewSethZtlgDR0+2kQ6gjE/aBvP7OABPW/MxFvkyoI/L/UIiHvDE9qXS0Vtxe0Tl
CKumHGEwUPziGB2UM095VWZObxrg9qQogy0ZpRTkBZsVePouut9Hz5uVmWqS1ziunWcvJYeeuvbl
A0oLPlRmUbczrih9FiNAw88Z7dCpvuafWc2MvrT1HhEWdds4z3EidejDUS0miRMFlc7aEinuec2P
FS2A+O+cW7kISU9VfPW2M4jw4IvpOH9/rSQKOBP8XgPcEZPWCJjTCa6rqjM6z6zLsFbguNXVtZR5
XwL9THT+e2jenomRQGkxmkI91WmToDtEn6UuLYKsXnB69kJAZXtCY6QfgJWe4+QQkUZCk4OFEwyN
atwJ9PVKn3+rHvt4Z+hHTk+t/nioRlSl0642sxn+BLF6UWQ+HjFqBbZmuM03i3aw1Zj1KVwjeoN1
dJ6aNAn6XTvnNAA8FNodPxKy7jTOXsqk/4/AemMnPRhioH63hcsyXC3pwE0uslq01OiRrqqKQwmR
4tovFv/6X2wG5Ust057OT4/9ALBTgsnYmnFTbMg3iMV4h7E/u5qOpt6pNclzaa9LdKY3VseVDmtC
bJcgZPqiKE8T+7AdIAZUgZInryFUQfmVEJKRqM/Vwf8fm/lQ5qfNmLWYoCv2MmvASEJ8k3xHVEmj
qy5c9w/Ui5OAMVhYvV38IuDNPm3DcBVe99+NRp92uzQ9E+wxkjrhRwAEaQiu/OEdPT0XR7UWEmN7
UpD/0uinXbwfTze2LdU2IxsZ6K/35DD9pE+JiB/IDsTeAxzwXvspkmj17Z4RK/RPiGYxB1RL4amP
GJFewuWZCkNZk6D0ODBcM3LAvBMa8tptXD8gMzYO110YUv/aP+9GcF/TiMbxmIHuqzDuBbo5zE8g
7PfL8YhRFM3Ad2u46K/1qn8e+sml5FDbVyOUiIxQTJJDqNyJWcM2mGDvd7QaUpzULPKbAsHdaxON
H/yvUpWG4+RIqR9J7kFowIa9QTQWj3xhRMo/eCodJXTjRcrYNhdeBAigFcm+3j9D9r1inbg0Rd1m
G1d1aNhNGUsmytnD8KRWf/5Rlr+x/hfODIX4V7NlCmzuVpkbT8IqTquXsb2AZrWgfTPtExLs16zt
/713mWE2LMpBHFH1H/n1SeW+0yiV8mP6KG8RjaIMMUfbhHn+1NlKhNKRufnIkOqfryR0qmbhTMZw
6IYuIRsVbSh+xMsDxnPL1WUKcvMXEw44rVNNE2gdeDEUS2WSXDm02buOo7Lw7rmu1QwexMU3Jzib
JRQrV95CoTPSp2wfcaq5pF/dOsapZpPYJ4RuXFezuKtrsvoc1xRNbLXwxP9Q9h9VUtqMfhES8KCL
C+jcTGGM5MMqmT0GAfhMxoBLrveFDctKu4bmZXfhkY8/he7qgSytJ8Q0O3EdM+slXujDDquRlbSh
juUaBFT8QbcTJwH3h9MscmNkq2yJNhGLexaQMUygslJlJKSknDfBj+sr2aICGYtmmqblxVa9YI3e
fIxJg21OgcwEdaZ0QaMwujkpCPMfuH9MVOv3MxHpmP0ZfCana0bVi0XV33KqVtcho0bCgMSOx8ky
7wdvz8T9RC2Mxp7N81B0YdbK4X7K3KjJ6JKOvVc2cP0yHNEHFEI2UzQDJn1N40eM731maQinz1e+
fds32f7gegQPbN1bJYJz9bAkZFlvO0Ib9CZipKaLiMEP18h8UkwbnfB50cTzm0wbXN0IylpCfLRF
A5wkDtbwdgfoQyU+EUBZ65rjV/8VBFzIipOEf6es4PMllRsp6eDYa1gAErosCGmCDIJ4RpLEFtJk
g3dH7GCmiy/tfkpxjqT+LBUVEyM3708zZDFFoJVwOqJOSsLLnixbvJGo0wrcPR7HSyv6aS5nVss8
RQ9nGdSp7rD+K+YbykuOWG0e/1tmIkIphkn6RxL89pJ5E2SwwOM89Ki32CEwqBqXeOx7+lKalPHj
7x3yil+AkWMPSIxpO2siLFrQ36CrRT28HQ5hu3rmLab3d0jzWqR7dkrnC1zDRA6aweUu3vOs6uc2
3HSHf8EBoWYHZwkNn7JJILETi4OMquZ19PfAwmuJznASWcfevxALJda7emL9w/DOPnSjEJJpVxRu
rQKkNzJldRBPDSL8DHBfTUQmrwYOQoRmDo2XbQiX2tmnMt4lln8TK4RWF1hhH4WMYR/q83qUMgLu
5nQywRfP+dOdkg2fSmw4nHoJT2gH3bilwShpRf6E798Vf+d+bPTLRRY/+m25spjLgnrK3YiJoJRk
EwLPTK/kjrgBwdXDm0KHtsuluDQ0Fk9MY28QN4ZGnTsHJ++I31qQ01LGURBp66LMTJGFdCh+qwJQ
XtaemU78CcFCoH482a4PzmoUWoWTCSt7+NLKa//c4Fz8KF8bgXmnVjvqUNUT0lYipVWeYjAbKlZY
eN4w7+VvIDyJGEnRxqGXoWMHtm79PdOZjhjdGwBLuo6SM11Iu1nluzCF+hQZcbHPgbEemanUmpts
1rUkVU7waT15bsDtEL0+Cl4F6lagv24v+D4QTpzlNpdfGS5iZDAoQs9uXfFf/0kjVZy22hHB/+T7
eSHJM2NfpDc3/CkjUxUIiriHi2yw3LaMjGi5kjv6BAAo3GgG2oGPN0l4CQsTfOIX/j5xenPmogQr
Aqr7H2uS2fzazGYMKoLHgpJCzPs9dmFO2wiMZ+9pxxO2FPU+ZW46ILwWmZRWgxmqaVRaPhHHgDOL
U6Acs+78WrLNDS2lrPcgU8Ao95G+34NJNvrzf9DgPR3RIxXrj4cxYgIZy85OtCxOjVAqwT+GJajI
CLOSSoOFodWAZFKaF8kUdkjUQ4nUOpNOgo00JtlavuXkme3MDLb44P1GKCLWi0U2wzYtkG+qEJnP
pse9fFgyjKpdclQLnHF6evS3cGIfviEvqcF3Lo/9rhhlnbG9qQ7jnw2UnqZwQCjAHh4mEJkXonU1
F7zSd7cUzWP+3MYv5xQkL59VLxxpN6QA5W4B9YUCverz42rub/IiipzVaDfFZ4h+9jraRex49eSb
wpkumYJi+TSmrguvkbip7vo14I6s/Eyx099FDcnFCq+F4csBatwhdJJkAA3iKxk7lljH+HLGQCg3
tz88tSRkbiepda7k3+H4VG2YsTCOZ+cd815LKTbQy2dfo6mcBcO6cPUbSjCJOERyiaHIU+8M9GMB
UOkKIlFN6+1jo84qvJhpTJ5W75NGeOrCliktIc7cz4EJRjCTGdbGDf3VMyETemJ0O2nQvvF/J4Ua
YneoeFL9a3xyJX+lFvNSlHyyvlTFZ1LTZvGz8rS35lYZYJqMI5V8TFZ/e3LMdOAm9wsWXOI2KqiJ
JCCbZPwo7f/QVGR36MxPvpZVeT++G81UooJZfSDPNv+LeeSAyLTCB7j6PiN8XB6GgIhlVeDWptaD
357HRmHX9yw7kFj1NgO4RvLYff50ANTqmSi7x0tafWP/pN0aL5oweeqXehHEX97akLBirTpoWv8T
jjqc807TtkYs0/WkDFzL0EJs3L3/9d5iohOR1JVLxBd2CmrcaairFoZOnKBFrr223n2AqKgRxs5R
jp253CTo1ijN5pKWkpruYIY+I5xu29Tva0ffY54Z/7EAFu69jeRgTZLZd/o2+aFX3Tjgk/arAOIH
FJmpgO534y2VEcivOKGf+9hDCru9WSPgJd2eaN9rzsMg6/dLX9X9woyto5nLm52Am+x6lQKtb5tL
9Dhh2H7I2MjJER2AWnTIvt4dG5OlzLvmutukJqSBjWpZUqFxzoj14qEZlbw4ylt6I1TIePN8DJeV
KLc8O0y+HRd88dlgxoJcuk57CGXcJnBuLF6PBccyZSTj0C+j3Ndn62M5QpX3Nxy+0+R2UV3I8KIn
KBDfKvKdHLbytakgN31/fWTOSF9V/zp561LFS1gvLOzhUxtF01y8lHxjadqeXm3PqGd1qKl1YvIJ
x665un0zvBOW8kYiQCGpUlqkbyDMUeQBV4300/C5/t1TnmMh3FpwDP/Ca2wTRwyShMdzqxzAgoX3
Bhz7rIqsWmxjR5UYj9nE9T8aUkSVOy5d7yaAI5CsSETyIiea/YymyXlodggFCnkqq1uAEbNBfgFP
Kpw6yaZrhkHgDlp3M9wmfpE3O1coQ7Qkj28ZSDYvM9kuk/rMCT7+fAA8wQfHhUmgLA2z8zfpBCND
SNKx3RKsBIL80HtpFyoqPvR0f/IagUcTMSW8l2N6kRJCJa2uaoPM2WVSRzTUDgiiXOF8UvygYRfg
EKv4r1SWBYxyLcqS5Dn+tViatsXmFvZjMgHp4AQvy9BJDduGLdY1LJblZtVsz3++CbHtq7WFiz1t
LtNhcmcwdHUsnzpmYAvPbAeP8uObPVZUkwlYzNsOa+B8YOx9hk/8Rpoc97H6xtXtm5FpY0oE1EoQ
B49RIqnBqMdjlOQrWrazQVd+c0x+f96ZUbiXrl1Bd8VJFY/PW3e+BvIFnPfec866EJAbJmfIYHm/
trOBREUowsmYBy9JAhEnQyFTPX8ykC1gABkMyyB5JsnNXz53yUaJ03lUy6GVgftH8ikhbaQPXT63
kjeGIRJoVX+eIYSfahpD3NbvdbHwk4Puj6TAsICb7QTITs4s17x+kY7hzYXEIKUHZ/4lPMBD0B1h
8aEJvZD0sMOB7c43Du0sO0F/T2/3cfAyeDLyfOZZMjuR4OTtmzbggYqSeqqTHXFoWJjgEATPIbDD
mPgra7xNoohg7SertLH17Jh5GIg1sLlVSBX/5bZyUpFeTaFFKdNBO8r0xTzlNUumZ0O0YS4t9PSx
YJMfeoxegu4my3A9FsvIaMWjXnIG8CMFxAAXiIVRTZKB5CZtoB6AMe5BmZN40JnprEb4ZGl1JEpe
3KFyx/ug/Ixqtn9LVQ20fHU72j/LMnJZ99A2YXrAt+vf/nc8gI4IgNBWohOlJQ+9vThdC8qn9rSl
peYPtfRicWVZksyeSZvycN9rsKJe/3xpOX5I/DLJb+w0h6OaKFlSL/RrwG+uF21mato9uaEw73h4
CGXLwdSWXXLW0NVlukYP7Qr6fUlA+6YS7RAhx2RoJhqkRTYKPVK0+OT7UzA9a3BNPL8+jCn1xSIb
EU7vpkOUT6uYIq8j+ptKe7ZVOqk1d0qUx6q/kIhwkgtslvb1NMPNhcR53rO5QpB4Ypf1cH6Ktw52
aMO4PpdtaxnwXEW3xREHmjB1Fm7Fj5imkYhqJqX1YllRk471rFzgoASpM1HmDmykDI2i0tSD2OIh
xjd4UNGed90s0VKmFql8DESlNILqvlrfyFBO1/B3i2nzSByjv7suxnxr2PIEvLTN2akwvQpw8GPP
82jVgYx4LuE4jCE18cMVXSNIWi1neuL0e4dTuleENIGjFkf359IoVY4eoIA07C3pasK46TPQiVgT
GozoIOoHWfMGaUMdHGgdKaI/sn3yveM0R4nZR1h8A2TCdoJ7y8c2x0an7gm3XsH/GX0SsOzEifAl
k8z8sdSDaOjYnHESrVIyZVraRykSmq3HYZpQwwun/WuUeJ48N5rC6bfC2aIH+OXWGlYnqdSCRlHq
RrBr0aqaLtSDVEUQgEIX48WrFhHWu6cT6P2ejdJ65ZDL9IWSnjMQyZcpThajqrwXoMUDGd7NtGGF
sS4euShP5/KbICQNDeqZOVS+PUbWIxUZNSOe/b10CnNP75Yaj7AtQDmEk8UPuylp9plW7xglqERj
nMGvPq+uJ0+mz040EjOd4c3EvW5Pi13wEqjDnvOoxyhohFH67gnc5SmpxL4yOJlb4UTWTz1SikqC
S6qvWFwhKV+q3UCMg9/lU6wQW4x/T/ffvOXqDwowLfYD8dvO5sTwkbfNy3sfnN5ktN/oRipH0Cfd
+diPLXv1IZwkMj6l9LeJBh2ylgLXZ1lQpx6CYvntS0mjDi3w2vmsZpYvg2ZinXytGwAx4I6SrIxr
d7IBYRnzTr/WpXqqid3g5XZ6B/YkB0BgkKNuRejtKAdJZtd/8G+vZjmA1Ph+mDpF/Et9kqQYmdZC
NCM5ULxxS87tr77EJEchRT+C4F7FR86KjRieX24nkjOo7P77iVAqmviiXSqBnK4uon1bbZSRQGHj
5ZIzEeYzNGEKWqlaFlMZmyvh57wyyV+sx5wNdYn0brSSbO034kr9NGx5ROu2uGDJfbgNH4FzgHXo
Wa4rTqFswU+KBoqBmeDxPfUMwiC+xI92iKU6xk+Zvhv/cStPPJuxa/heHz9nJcDctmh4Sio0IpxS
sxEmLJGZ/4DVG5ipzJTBjWa20F3I+nB6w8GhLjhLYUbLmfswKEMAV1q+RXPUza6hTlx8UBh7FkbG
/sVaKJLroQUuuGFus05E/8DESvtgZ3ZU0HQLAsGyl4/AsihbUj5K+XxXlqT+6xUlzN7XmrZohnM4
3Mx6LCdZRUluXI29bKcOUBoindrFXcaNdZ4qGt4VzEqxuQcF2H/9TK1OW769zgxoGa+bhhXAFBEB
PbP8pcoXPN6N+Q0QsXTPAXjAoD4Js3OPYVvSSd47LkNvYgQBFDjInqANetulxlZewgA7rdjLGs5L
OBLDr70ujVENYTk1tYTgp1nsY+b0Mzu56hZ6ZA15lfrDybxvm3YF3Hn+9pBu3hrdYbCz2YiYmaGp
nPTAI39snBOYHz/BQHEt/RaAYE5vwn8AK8cQdrJTPgdn968EBiL6bMbz3puLi2ta6IMh7STT/SdX
mAzPxxOlwrEG9Y3z1ZozuHuqieHOo2570q5E33562aU0zu7URkLnZ/ZgkjL2n0Ahc1C01D3ouSnS
Tq3a6q813qBAMSbAzUdSq6gEhNoO4g8N9aSAUQVPLT4AKdTUSRtdgnvs72XYSsWXQKMKWR/mVD0X
SrtMLliE92xKaD7a4pe/z1tGzD6r4/i17wPfSvcJSWVl8pRcQhHXBo6gXntSWYgFmvupfV0hG0zP
/3aWx4Poxk0YfUwtpdIVpkPsaSCzX0xNkFE176unYKw/qg0iXTQe20qb6hcQfGlb5J7qXugV6GL5
7zCvq8evcHEBSrYtzKkFrcgdo7rQT5eZM3yr0lSKyQzDjDFhMOlQhln8Hs5Pvvrvb4oOPDlkeR0i
CT10Cfb+/mkVZM+RVA0/Fxl9t4RGh+3e2Bsc+b1vkEv0Bv4UYA+2vl7Vw4KnGnUQUFtsFpbzofwi
3inDTwTCIhl6O2U0jVve4zE1MSQNl18aW++FpZ61nIPbfFKPYN55GLw3URX314wKGWTcmi/petFU
2OmyoOJ28kdzgNBRvEARVht9lu2AAfvyDY0jCv6Rupuxz56Yw5mWHC5L6nnxCKNvSDRQpaY0zrHp
jtxxTg5NJsJA0KeNWT7o09BsO3ZeWlr7TIKg3bbQYgfMRYvgyyUxSos5iJUotaEiu8OWq6j3pZr1
MA33SbjPr5GoDr0Eb3TDsPfcQXOAkzGF8MCROsbcocOa6Z6b1TT9FCMFDWrNGQHZreSOiBpeGoKb
qrgtpoV7Gh/sLBQMJx8tbKt773/yJREopw98tV5/FlLOYwzzv6qnRGuLXjXjtpjq4+ZjoGTFJHnc
rTRhy7hmxltnDOvnE0e613MOozZLjqGqFo0g6N5kxQzReYDQIc2f5XNjmEuUrb+JJ8GjMvtO/ENg
NQwlPnRcY5l+mNzasDavUVp33XJk/DT15ffsX5cRnL93yNnx6TxTpeWC4Mq3bOg4bA8Wl093vNUX
XQaw1KFmrqZDAfRW1rnCY8/8i17+gOAERsID66yctdvfxnLg+NfXbasrz7AVG4RFY1KrQcg6JHBM
Rmvr0TLfFaw1dUhO3LqcuudxxHPZgIKNzWm4FUmixt8izW6oREL4nRc9GCXawrsgDbMv1Xf4kElY
1z11UFdWirBsdAwjpkNOcLuRsNOowoWum6QN4sp7CLr5mfFGp9gPXV5lPGlywKOCVs/+SYOIuSmy
SYSJzUqNwDtPJAVvpmGzg1VjghTwQ7+Ys/fIk437nO/xJqLadS4x37NSDjbS4aHfe8fFeNDbCf8A
QOheuSbk+0W2IOSHfkzx/nSzo3+BhsfvupW7eDeaD/Koh0U/Qy6/3fAoGJdinT+GDNO2JRsxaSuH
fJOECe1fHnoLsmrX9uPMgNWMRE+SIp5PsKPfFmKK9DiaPf8wcjKC9s45mUD2c3dh6f7P4UASjwva
TyoMjJcyfFhw/Q768ldkP9R+ZROOPBQ2U1oLBlt2iqcmBsQmZfXJLhK6EpZPESORQc6/yqwx4TyH
Il3A8H1kprlowpUuOmgRoxpcwZ7TbMNnaaOPMUfw+UXvUnS3e0uwKtKIq2P5hdkbF47Mmh97jYL/
OXKd+roMuLtLplsVRT94+E9pLScLXwFpL9CIZIRyadtHYcX+NpogwNiHnPnht2SmPrbFwTzRVegX
LTq/7GKytX472T2WakDENPwKSQ0ztDiGVrvBsibQaaawre6MjdF9vrScdPeIr22M7cW+dgMAzvup
zOXCfiJLyxdbQk4jwyY3N2w3iqbo0SGvqC1YTbYIanES6T4uI5tRiFCiJy/XeXxTl+kr51HuPtXe
FZ+WVqxSVUJjR8+sW5vo5e6OUZU4RNBu1KgblKhlImKHipApv3YlNji5w6/etgUNseFqwkBg2faW
2Qw1kgoJZcZwnvR3JpEi5jVzskgyuERgcC4HNONkfWTcvHchxgXBoTeZBs0+J2djGcKGOcqGEbUa
vUV2bxUAO1raGbsC4mi1BJnK2kvJIle4Lrd00jpKm86/EyAzGMn16zpLFGV1Hj5TGA8Igm9MBxj5
VfRXM60sb8gKHS1glmwRKoY1QeD80L1QbHelXJEdfH61+O//5QX3vwwglBjEusrFArsuZMJZlrhN
0tdV+srNeGlALvBhFwpAlHv6UaarkEiXaSldqfPGfz7AccXsaha7PjPJULitd/l50L0BzITr7eij
a0s3PTrD+5ubD/gcVsKgz6AdPSl+HSNNOeq1i+SBMj7sS9YHP3CHcn0sICxmfTOHwxKWzEPRj/x8
fu/a34bEOZ/OICYu5kzlg10a7HOwvDJ0gUoBNrBIlfiwOyIjBquFR13KE59lgjgQ04wOULNFMo1e
ACqktU46VEuBRTQuZ+9+73UEoMXEuwXt0GZBayBOfoZT7P7OlXiedWsSLjVCZrqcbVzyWWbDdNo4
tEVfhQOPW4QYxwFnmNTdmT+X6OjqwujLYXp/+42zErFyI7NJQAhULdVJohlYbBOLbfuteenzu7Zc
V1f6S+2c89rImRzAhqzzWJ1LgfAdder3OlI1MgDQ4lZTOs0JInvr+wC5ys8m2rUcCyzePnsLsgIu
oa1+JED8KjKU16jWaYMu7ont+qLJYOrmO6Ys6ogTuXsrN7VXNyzwDy0mHy3yI8/y79CB9baWdg6x
N2i9DidcgySXDAe4Foq3RdCVZb7+I3ryiSPVA0KdAaaUOj4urEbsCb+Q22jJ1ffo8MwwAPaBL/xE
q4c1N8m0qxoXYTIh8axLiAW9REOVxCHKJmwJo7y3Hn/NVg2Uwm7zrHc7Fg28Y2w6dR6o1yQeIQar
1Wz0Y/QPEhRzReRJW4hIaLHB+W3LftbE4baIoRRW8rAdE8RRAKZ0tx2fhBBKd3FhosR8utPqv4Cq
uWWcRo5v2VQw8XR8XXAX6CxBwuh7bUBObA+zj2zfWoPc9G2go/mkeekoPcM5o0D2ktjbjvkJnWZl
JDLUVMiKcbgUB9lXSuuqjphAak2zf8IcPdYj0SIs4fYCMpBA09k8eC+JLATcj3KZu+KuH4rK5+cj
FnxgOO1jTj/1aj/0xPVgXsbJmjVlg0sXJNo1dTV4DnXPMLxEALOFyhVdCIxkeH/rbSQwU/Ir1x02
Ze3My635D9N6zXL2SYX25aMUycd9o/kInRU24ahztZv8PSpFAkpega7e6lsmZ+/YNqnkGBew/N8c
xF2KJzRtn96q+GMzfJ34v7gwaDgrotV4+gTtlCyg+w6utbpTV66a713XX14pdzfa1R8g68qJ6p2a
YSS/5ipRBpiVYEf/m1hQ+aFVGAhdLg00Wy4AGzR3l7P9NAK/D1BL2bBDELoO8W5R1hFNsmzVI4dT
0LSHP8z2OhElLASjf2Y9sejkl1mGSMvBPmEIcyyTnGnm7XTWYDA544KH75ufeASKBGib6sqvojMa
Ajx/bYpHxd4UKHFjJY8ikXS7aMEz2/BM2ACrsW3me5wD3k7bbaKxGZf/Y57udSjOe0cBWYY39TE9
dUpBI7Dxf3go6v0l3E4jX4mybheQloJucXhAPpO6HkQotXRDmiiPWvqGVTXfHuR22pgO7nDSMoTW
yFkMNX36Hsj5YtzGzUgxzdiaeRUYQVTcYk1X6NGuyBGafzICAht+HmY/pUU9okSDW0eFfMJ/dS8b
O2f8pouUV/Xyne820bohDlbcUUQ5NNSYConEHx2AyxSI3Kx0kmpW33moBy9XgaOaYSSk4OBu7t/o
nrEiV4znLoVdO9kiexR4pVG/uv6tvtUgsxigh4P/WSnoshT3BLXpq/gHco68AlYemA7UpyH4YiRA
oONkiq77xygT0F1dHkexV8skEC4sWlJUWF/nbxoJrYI/IJQaS/yfKSXjLis/mveLQuCOvLkMhTvU
+l0v/vLw80d07o7qPH68dgBubM/u4YtuUDAB9cpIqk3EvSqZnY/BHnDYgrVA2nzt3KOHcfnYs+RD
kdUOQRX6jHZD1Mm03X4WpLur6YeUFT9zotQlwSmgBi/3Er5VwSc0w3EdmwzOD9unSNyJaSRu9DNH
93uWNANNFj/amlySWfqwRyiSCyjeQuhSwDvGY08iz8Dx7yFEl7UjLxfRDJg4ldFp2KYMln1vQMuF
TqAR18BLnkqAevcK+BaSHd+2jxvs3aADoxWOW31GIqqoCNMvBYf5w6OKvMLYbq1q2T/mB4Ss3EUZ
QHB2ed7J8CA591/vrXSMZhLusXpNjaSD0/joHuPt6rfrI6xV31t/frPkOvwKfGoxv5HvQSaf8HpD
BpIryc2hnvD8VbaQT+kmMRZNRv9KFrz1UsPpae9LSOSzPEGc9gUCcautuUl2ufqOhSskYmorlMX/
u5zCeQQ2+3pm1umU9PoMWfCZF7IWIKiHJdeIyoF/+YH2M1orUWMACJQlCUdoBYSNA50tZzxGFJtH
Al8ep0xKPSkVnP2MrlVmnnH8E6FfHVeFRlzdZ3EhnbJiZxVfezpbwCIEFTP53a5TtmRFfep56P1I
9mX+JD14Hypy+ixWD79fqlt7RxQpeaUFjp1+kYi/8hlVsYATscofs9S5M/5xxGp9XKK0O3hJKgmS
l1gPtatbTUAnl+wtgIaicKTnNA9BCSVKSuEg9I7y8RL4DMUwmDl79rFTeOv+3FLAFMI0HsA6v44c
M+JMS9W0SoU71m3TMICFSBhZK7QLKbt2hmxvtwpLZXiT6UNIZ5tvUOMWfqu0ftvYbFnPpU37NhLl
QhoiP9YTzZpcc6VSGFPDbcc/KDMoJfgvAswUU9FkAgnY71xUbfqwZ5Ljdxa9yGcGAmPW4N7Nwbnj
E70H06emSK9uDQXXPboOISyMP94OjKQ7R62kp69E5SF8H3P+4gQ25/EXfGKxbz9DdgMYQ5ms0dLw
7b9M1pet1HRRniFf8jGPoHVzdwn3lKI/6jz699aVMH9nA9dQGyBNIhjciidsSMmPHLE0Ytcu9N31
F9xh7foID6JgUZyED1eN7Wd4T9KJhli/mOGldwccHAwYOy4y4y+8wika/2PkvtRi47ccfQ2p+BWc
SEYvi2nLS1LPbE8PzBm5iuvZRyrSepw5DW11Xyj4WXaYf9Es904ORX9cEhcuyRw/QARQUnbV7mO2
mFR71/7Xjox6Svbiwvpo6OyBGg0mKVaEN95eUWV78EKwxzB6NtIhJFODgH/ep7y8LneVh1nsBXDl
E3QXnod/Sfn5QDa7MPePSofY3Ro4u2qmYTLahJwBogVVZZu8IKsCUunqxyyuJn+yFVbte+BcwaUJ
boramIu18v+HftoX/iFBa2zvQ3MFroSMNVSNepdUfeIWRNBDn37/kT9P41zWxAsOfPOqQvxVuzX7
72ck+lgxDXtgXkJrlnVMOLNRF9Q1XVE0DkQxqMwma7qfHBC3LS9eKNEYk7QybfNhdA47bhLrVZCl
mdbVf6sW9S3qSsEnqkG6nsORZz7J68AXGuOJjX/TdmvxdEWFeUNNmCbDI4mM7sWZeNyF6pr6Q7nl
5euv9zB2l83LsgzyuV49fG9ZJMknJQnnbTQ39I6WcGY7xejZAUYtbtYfmI7tF3KjPOyXwqP7sVun
w0HSuuFJpzlj9f1IUMea9JNmi7rMhv4MvERf4Vg/oo2alhYkMsOLWLu1BEAEr3a1xjF869Bgeb0/
3GObOt8cEJxbqg3G/nuoKufyP0XVfgM/hFWKsJ1sa94MlPJHy5ySvxv9QkG46vwxttnV9oarH7GK
4zmG+TZ0iolgKkHkWzfreHfZ4lpc7zzSNdZh196E0i+NRm6VbwiezZ6/bhq9GV8GJTxm4Orn1DcU
6KbZxQTk8qJ7wBxK3WszU2Xc2+rX8qY3PV1j/KW8yPXns+tegCtP7j+p9FY6oMThfrXGVfI7dLYA
U0YRoXNvm49D1Y0//cWebZ5GCF/L6qgp2AFmXcesLBBzK8IJCRz6ecSImHNUZQAxbdi2eq/lGHWC
EBiFVmaAySgLSPRlIOWn/QidgE9WXQ0v5YZBA3SzSiz7DhojL6o5mzj6lhkxvLwiOwYY2w1TTkxs
iEKe9/Us3k4W2URzFv6KVyuk1+Gk0IXU/j8gdRok251GI3iKY6ftEiDGroAAJnpM7UTXkey1x1Ge
j6CgRN9cWslhkq+tKqTtejaq3SiQkmTBdNIbb7M22kGBaalPRKxvtxLzScaYLM3uBRud5uFGLT2U
XqJn+QQ7ZtaHaFjl6uixNDJpJyZSU+ozfPRMT63eshr5kE6y8GSEFhrGPvlouxw+/DMM4r8DNRDh
xsBl4bmr/HnlpIiDe+sZIQ/xtC4CqQ0U6C0cmho8M4XunhztN8ypJhKv/BohsndGOIyemF7cNPKr
V0oJ6GuMi7fGI97etV1HjyZ9dwabcojaOiQW8BEYvgPWjmh/AcuqtJH4QVIo1zrpU8PIt58B5mgX
Gi2KBILT7bicNg19VsUk/eU2iHE1lYmEkE5eaRRSqhj2L8MpZCzUPlTylppKj/pxkvHFNkh9DPTU
Y6KzPo8Cwebq+ukwf+8CrdJf5sZXOR7tDgFfFdMSWGiUkGUos4Hr7Ub++jbMGyXliTeUywBO2VVA
d1TMfwFQp8mZinxP+bPK+5Z0PEU5GXA233z23kooYORDPcHy0dYXNkXZs1/y9t1t6C+6OdiGo2SQ
razq9F7yKPT9xy3fb6TzcI+CgaFgq8CxeN/t/iia0MvVGE/BB10x/hR5ytBg32gQy9lJwzkbcxu/
lNAHcMj1WYgx0phE1w4XM2ggx4ofsRy+zVLJ7BUJ+fIOzoBYfJheFmYDPjlRvwVWK6jv0wUWcLMW
/N1phaqs4PDObQwecok5xMMX4TsybDXAZkEJtOx4zrz+vDx39ft8Ojdh5B+pxMe8q8U3pwLn4n1j
vO4LWB5tb5+4Mq9jrZ+wKMQe7OKJk6pKWjUFkS6uF7jWPzvPCCVWxP7B49H1UZ0E8TRMw2veB1t8
R9NnYSWNMkFuA+LNa8iimCHlMnMqM9IJyKcq33Jn1Py2TChKOfgvf7nFkNrL+OtUid2Ns8FHR+B5
4DWpW25mVkmvKYlmzTLbsWzyw0NTacUqVokFAIsCt8JD6qGQAPnfgcN210K9EXLfbWxl8WZTpJ01
w3MHF7PK9N9996tgndamy887iL3ymeqi9ArL7A1tf7s2hrmh8cORQBYP8EB+mDS+RS+BPxATjwIp
GmkSSmiAAR+xf0sbxqs2ISm6N98adOr9KZvSG3R4n0BmgQZIi5MLau4RiYbeCoCM9K6tasZ3F9TA
sy4hWb8moCECVu9vp8eBPr98jG/Uyv9o0Os9zSXEPmVG5T1ecgY7tbSX5Cqy/1d+8xeP7p2sMrzX
fFHRNN9XQDF33aRiQUy08ryeYdSHCPCOi4H8z0dDFWixQisKl0WJsvkCIN+ettc6lLm84ysFmayB
kQi3HQQPO1Tu6gSu8TuRJ3o3Pq5DugVbLagmP+gME24Q6x09CBL9gUX3vlnJpYv8t/ICA+ylYmID
eAGqgGyDXHEsGQME1i8RB5XiNKy+9S8QdIDlgnrcs3SQNmdStJvPuPq76zD/OaHeNQs1z9VULWHP
+ogBmsgpyjIi7jKZ/MD7njMRdbdw0svYQ9tdO/Ss/hyNmpqI7N7DkazwAFJsJJzyM8t5GXlHjLVa
OYOhF9rWHFEEgQvmaEk+1dJ4n5ybpks8aJqVxWbcA38rnS1C5FJIKOdHNn2KjcT/JYtQQGX/ZTyY
thZx4hYk/JY1C/+cvdWRCCZv9gn4TDwZfF0ZgrlD14xen5Gt3aQ1vwFmW2cb2x2deY0GSngBPiv0
cRu5UOsbGV1c/MfLPV9GYZblkl4V93nc6aBSGk745EBZ8QLUYJYmGXHqJYA7WDst14DG2frILwmN
qPQKeaEVcK/+ee6/v9oZXzh1tSPA9cPcT4t91c/TVYgBGnKIfWqXlBzun4i8Xbaq4ccGQ+5Mt1YM
LdRKd4lWTo99GfwNVH4h8GPxwEdobKSSFapsmZSo81wvBrU2tdIpcWEwGfe6mFeL/QlkGQazGt94
vnEvcAL8DX64nBgJHC7w370PDXfMtiE+fzZfOKZuJV3Sd79pxR7410+yg3epECFdtxWoICtehH7n
56vpcOEdEk/wlbESTsXpXgNlm7E6szaFh2eC0tStJS4bQZWYQBIpGFAgGMrRVsWlEkxXcXq2ntMl
tAsNEgNvZ2DbOoiUrHpaGm4CRfSSEtfQIsD+Yq5GoDTtuo1FFJQYKgRz48Ejo66HxtBg2TMZAceg
p+EPEgbAbX/Kr8dhy3s1XTlc0WemviSl2lCUxEBnUhajXrACzbdvX/rHHA4rftrNZu8hkBUEUTt/
jLafX41tzhmqMm56ywi2w74iLr4ZNzjo2n+KBdcHWSZgHVHmc8wRBZ7J+uZ+CtLHoRB6ApV8thUh
xQEhAc+Z89GToz9Pg30f9nFL+3db8/yqut4POXqK7SfZcWLj6gSk5/SEoSGmtM3cIZCppB5Vbn29
DgUzCcC9DPNyrN5qGp6I4k9CBuAw9Ag6g/BFqNf2mMKmvSf/TohgzlJPg1ah7ADHRms46x0qdBSm
PqbxGb8y4WnlCkqbMGhibGRe5gKg8ndIwuTlBc4IYgfLAgQHKms/JPSiubP4UrMBv228jsvpwNie
2wIwRm9pvxLC/jbU0l+sQkogF2F0F3/Rj9hjwMHJjJYoiez74WoYhkBI+yJJWdfnzqYrcJGWjKyw
CaigiSvKEpvA7zmGfoGKk80Ni/tfDWYwVUKcZmbr1beRqpl2LlR+l5ess+YRn3E/KQSTRvhje/GE
wpZRYXTk6eoWW9elDtEidU00P7QRE7ZEVan3+l6VcqAJNa/sV0Hvuiu/0Gt7WvNFnwd8Bq/p9lEz
UFiO3dmrCXpOrAN0qnDk8HeYatQFXvrEYY6cVobilQazGqT1kM83hPoLf9bEqaMS0FaUkm4gWfVD
ltf54l9ObUHz/ZvxmYoRSSMT5TbnjJxnj766fFbqNtbbNuKQWO+tyJCm4KOyYIo6/7tkDiUfg07E
gVbiZ0+vt3y7F4wV3+cwD2z+S4NhUKofPNNATb3gCh4vqSBq3zmrhPbIptBpMLB/NDHMrnmh3sZa
SVWw6h1dF00dSWi8191DJyI+2AkQLdExpis6MaAsadzIMZdal6NGeE4mqK5HjfmYyHintqNNPc0a
Dmt0xwcLv4z1YHbuA6UBunTDGac9CRBPBa1BkR2XdZzHinUbd1tR49/4fkmaEiI8pghG4nacPBNo
9B/sE8h2sFn2emulb0xvDGyTK771Pw++14on6e3SDfDLb6Mdo6joPqhXXWSZEcFCS+jAj9NHng6a
ZiUWtJwxv2/5oCsIyqPSFce2zfTJ3SKY4+hoRFdj4YscgXKZoGYXCL/PJ62ohbXUX/57orx3pSr1
ldUCJNpmzVoEWGEvDaEi7Mv7jg/cJtT62aPueh8+jUELqNJj+n8AIMHBMCrmlpveTR5culD1A3R0
PaSYkanOgSYlyQ0WrGpJ66siCsDK9W2AuAhZEiNqCDR0FQGMvJH10yXcjeFLDPskWlGfsCBKHvED
9myAT4XVmAy335ADYOZ0/K8EEq6ryFfcx2oCtecmU8ebrcgcSEkJwtMNkS08T3hd96e3p/P11NPJ
28zWjxvLgxjoHwZ7INauXQuecS10GnVOaMHdPBnRL2h1Nga+Ra2rFGMCFbvPc289qCtHimYsqGyL
6QkY5Q63VPfObwXG5RQj1dmy/v7yH+t7dXA/FZom72IZnoDjIQ2Q0K0DM3LSgH9L92sHnqRQJ2YC
tbleS1civi912WEvfOEAnb3iPLAh+pCyV9DY8Sno/J2EeyJMLmWIgRI+uxNVD2nBwurFh/jdNIMY
pf+we8TbXBMbpJReA8zAWEHeWRb8+v4wk3mPA38+eee/fmuL+DefgKv9XVSQcNqLMFBMza2xvHsH
oDGMW89fR8fkkXkmkMEXS06KaXWPr/tLJsV9wl7ZcIjzA1PYqfgq/kYdowHHudjtSrQwWrqWUrK1
aOcBdQs5wmtJ2fmWVBCDGq/pF926qyTkFLegvmmq4eiVk35lKHSCM61l+9mpGOpJIAY1kKQO/OPZ
814aSNlNrJtFT39pkw1x2H1YqBk+LZuQV02CzXnj5dZe2pq0J3H1tjQFhsaE4XS9yiGqhP3uc1Wx
rfxD15ovvSnPzER6IpIhKjeZ98IAMmySga7xmKKq0tTb3jOLvGJWYHCWnSffc4/ZwsrzhV1vy1mA
SFyEsawBgjO9LogXHVkjKeR+EiHFMSmfYYGIqZthHqbN3d2EONoL/WB5F1ffJ6qDJkTz/eGpfcq/
A7+E/HUG6uGv9Q4LBPjDf4czsM39WPm284WwViXwVnJRcrssUoAZS1f9cvQJufs5FYhl+f+3G/L1
2xrECUhmK4S9EBHYyoQoGkSSc2/YXNsO65aM3N70tocQYuIl8p3if+cqT8CN7gs8NKTtPGmpLZc2
mFGJ0Z1cttvu9T/zhZ588R3AAtANXqZAm53CQTukUQ4+kNXaD7VxGPcCa4rmsoAV4+MGldtOVaAz
KDlrv6Ssvp1NxKn0y9rocQ7dtJJwKbL1OKFM+QAXBt0SH0tMhItYLzqZcSwMFL+Jvklc3wCobKnW
PnCT9nWAmR9/K1lyEtPFaulvFkv8JTJFDU8i0GSM+mIzKxb5+mFCJ7BDAPgDseVkx3muRO6OFqA+
M3s8KoKd15RycHFTlA4BTUVOqn54r/ub2Zg3oqes/JE0hzQoeTjOAVF8zntL+jpleMzsl2h/9CvV
YLNVk7KDqK+LEkUtXXLIhIWjxvTsTGihg9oa5LhVct6uKbmk/TueIVqK2PQFM5gtLteukB/pfRsH
Xgc18OpCg9Teezq/yi9dugpJX9QUqRUpZM2JwRmQy1WUKqreAQysZlRd7UQ58XvJIi36q/b9BiiQ
ckX5usaIyD9g2t10HYczAvqH+R7Ze6CoNu1cIYxBMX3lfR0987YBdBEk+CPGe09iRcwnoSM0Mf2A
30qd1b82jEqbwqrDEXa7IjXLW1NYruTPLGLXQWSaSytu18QNA8oQPrmoEn9z8aPPOvnMUSDykJED
JJ+I4I4LX26XzS7EDjcviBXj+Ph922cuRLSyaazlxZOUnooqMfjUKGfFJh5RYpiz1RplVPB3W3qP
YE8cRNpMeEIa70VPGfp1BtbQ9oMb6njBI0xgE1EyNS2Tj8QXyJXqL9shbmnfz5oCpqajPGqzww9y
qgxkQLgqRy4xqamOe4/WxsPyir+NWj1AwXGi4/oozBZOe16jFiMa2Ea3MObLKHFGAnPpGpNB4jmd
vGbyVSfKXfxMcRE3PFxJJ2X8Ho6XF3alyGIB0KANX2RlCRE+zWimn546vHkxDSZDTQzen28OQO1y
XSvgk0f149WlIr1MxmZnfEh4hzgrxFIUdiQb5oUAIEdL6M9nqlOTCKGGE+pPrjTI2Jt+2d1yz61D
iR4uewASzG3MurPDYIUn0cch38ud3ZWC50j2Gk5pApTXj5js1oJwUrjTN+/edlxpg9H9nUdj3Bd7
k/a0GLI4r3Jz3VhW69ojEzlsD0b+vqVo0UnkAbz3oHOUjlTqC91YyMTNppWww21F44kULkZZxAvH
0eZVtWj6Iaj/eoWz9bGh4UXCp9EQ03pOdW9IlKZj7cnbOPNIbYUCXcAKU6zSHm4bvbMBp2kHIRy5
S5wPCoLQUk/0DDHgqcWojO4xVYKVUnz0RgPZB3S9zUn+ggBRlpjDy6wkRcpg+Xyx6l+YO+fXZ3Le
93eJ8GRKw/Dcn1pC34j0I1RQBWEokrv+yU7PRnzu+GIJP5K3r+L9tj3GM6jZ0tmbNUOkPNKkQpDC
ehQ1556dCMWCgHEqw4+eRq2Jf+zAzs8iKh38XjEclIC5il1cStcWs/yrNkeH2lxo+VecVDbk3aZe
x9ybJziUVagsA28ktFB+KqaPWhK1p6qBqTwFPl6+i0A5dMTSLLtqx2UBwXzbio6gSB2BPDr9fL9X
u3N4AX9dHcomrM9FXtRpppbe+6wCV0bDyYxjm2bVHWj8LyP31+KxZuFZLvabz6X25QFuLtAt2hNg
nf3jKFe7z2xSZzNZSbJ4WqGorJ3EqHI2t1Fd1bVn3CXd5sCa1ct6yABjScDazIdtqHnCXtHeyytN
R6SDVUPOnLMQSeCacAneOfSfSBfSmxxNfh9rzZRK2ZrPkxceUIbQ7hTGTmvco+2HjvVzmZuhOjQv
q5vp7o11+4+yyNVmIPJQC18vS/MjEVParDQNsm+vOO+TXiilSFyNQOmYniVNK9MX5qYpG4MyTsAg
wLDHEShbi5FaPoyCli/E+xN2XyIVSSniyWZxbi4X4lsecMHwIOxY8j3vWuqSB0dV0eoP2/sAzvV9
HKSSa0QJ0GgOu8N8/MfdTsQXKby6egZ/G1LGJ6XJ5pCrwRvsPW2IXFKyrXQlyRrgxOWMr4gOz9m7
VQ0PkCOdqil7XK2GRsxfxCK8Z8Ps0kvU7qL1Szm+pUOTKNP1EXjuIbApyMf6R7dfZNar5gAJz87J
AdUwWgVs80Z2kXU0G8ETv+bNSbam3nboLjNL6ODSKqahV4WgKEzajIJf8R1HNVCQ8h6E9EaRrTY7
QpDk5IzZ3iXFBq3jFECVU4wsHMubC9cxfpT6CqV3Jptl+rak71sg06iK/ZShSqr4geEw81CBJ4eO
Z+ZgLG3cA2F8qbj3HKOVsLnDicEsZPhevnySBO0mmqZZrbOKfkFhc2g75aLYERhJCQqw5muhEq7p
1FznHbxddZ4lHxJ/suy+NoAyapJQmGza17LvO4WvPFpHngU/5hPh/FLIMs74W6EfMoUwvEeoeYr8
tXd6iE4Us4Y/gQ8ephg0RhmFQdqzuFK9QMQWhYDpCPxas4hlHpNaqkGiVtzrYSqngEvL25D2JT59
hjgMXe6nR2hp1BJsGMmU89Hq5vdT4VtQqCelh/Ug9kzwusaEGKKRArFgw2wQJrJjauU5E2RbB2EQ
Rl7duMZZpnN9qn9NuKfPVbYrt5ObNhDsUQgmSaR9kiv1BHbmZDjvQXCnKkaHk31I0oESB/vLM84y
KqcqsHM6moyTyosSYCsIv5bOjmR8pOdk8XyMWyItXYo0CkU2ECwE+h2zJF1wmDGEkTYVwuBgQ1D3
GQ4dO2WEHXAicfNzP02yp1LykoLXEtizk0wuOpXAQ127JwF9wpPw1REFYLvSMvxVbXq7wtjx+upi
M+2Q7GMdXeme4L0bl1tHH+q96hkb4QJBuRLRL1PYdHyLm/UOs11ffi9WOsxE1M09PK6K3mvHw7mU
MA4kcroStuamNjCxvbRcr2dN5+0JpIGjU4c5MWx0fIgrD6XGagvqVL1uCLTpt88kFIJr+InmXSny
0D4SRmCCG1XHVmGPRRYLrOp6xlgueDIMnMlRqg0kl1+qnOB2D208Zi24wiaceZ+zAAlzKNqG9dya
s1fNydpAEUiXG3m3hr7LdfQV0l+rCC85gLhNOxoG5XkRhPDiZ066Xx3ctV4cwrDbJuyjahiWGLc6
XkpMwvZh2iqFuQlnmtBxXwM0TMdF+9w67O/D7teouWAdeH+oWCcpRLm6bZnatntxjcLhF/XFYfX8
YnPWKLWd+l31ytFnxCqVrzkhpbGAkXGCrBHBeH/byp9kodH+V/zPI0HWLKVi8lwBUP8Umc/0Xw+p
0Lm/Tk7gbzZPG3cbFxXlxSyHUa8r3ToMAngsEq5fGRsCrq+mYWBrKG4jTjdaDTej2O1NqBD+C8f+
/YEuAzWUd+yM1UsWE1yIh6nPzJBWZrY9wPiekNute8Uv+7AQzRrsJQUWsEK++56EuS9bD2P6zu+F
u2ltg60C1CxV39vzhZ3qjjLpg5qs+7/NIf9rVMpa8JOuCPNsIU2TecUpt1RlRKYEafcAJb8RwiHB
RCb0jsRId4mrEaIDuKL8oayj9Yv6sHEYC4Ttk+u5jdACV1uoTPJ0dUzJfi6TSim/cC0jmqu9/db6
5hmPawJDsz+fgi7miQ6HOQo4aAtNMyQjjbwMgvp5Ig4Vr8XpWvOfJQ7xMrtZKNK/A1C/uP185FaX
JRbfzjSsPOadowdiFpuUILBgBJggCZUUT0BYNT0TC0zZh+P/8R+F3Q2+ATYEbnW+uPNJnbov3sRn
C7WfIniujmN3YlygSfHrAyc96kbRbaizVgH6cvW+DETnS+xmPGDbQ8Wrv2oA1RALFaczmRUwneYE
kqkgQ5NNS0Hjyw29u7vhihPdVckYYy3cS6F1PdL58fq8bVsepHRMjAIKy0tUQqUIDZ71BKfjziu/
87xO7A55xqUI7QHnYdrFU+8RGY1HvUTiGvGoCIKEyL7rNUBPYZYyFf09s+Ofe9YwnKfR0Nk4mV46
vvjFqRWVejX1lhipbegmC872empVd1FyN0iDyodIcyWMGUhXRp0PaajpPBP8+Y3UzTMcBV9vDX5p
T2KHFDCIMOeWuXKazLJcYbVNQTCLS9Oos2/rheFi9QkhoTxf3uaKYVXrcbZCcAsN9QwTK44fhBG3
kQl60jVKKvGpY/nym7pfpT1Hu8WOg2rXOoMbh2N0BmPMarZQhKDg3C57yk0WFl5xWG7yzi7sQ49o
5hnjNxAjIEbwWooFDOnPrNMxKKkmGu5jIm8WviJ83lIPU3ZU+04wVz3YfrDDL8oTpMy4dF3e9zzw
/gEVcAuAL0jNt8bGJkMX+Bn2W20lGf6d0wuepwMH7pMUpNFPhoAHA834qgbpHop84l7xpg4mtx2K
bZQ1BvjzJLbfyyy7XWw2xlAGPKsPM5Vn1k57P5V1+7GPdpwqRaQt3YkHPCMmya9WfhDUuKXr2tVi
X5f6DNGYtEHKrYPjaEGKQuIWOD+QG6DTtNNIyxd18I4TTO3V8QZ3Vra5kyb6LYRDin36ftxJoSDN
GLA1Gz1L+IxQO17b73r6xYSBNKFpxMrIaLs6Jfspe07pon5sBn5G8cvna59BLORStx4SUT0ALOQ5
7rRabwRfWQ8Q6th4ZRJ3MClPkWVf22oQl36twltZahH87cJo5HxIOxuoDD0VVlS2yDtFf4gkARkT
+EXmVkbNwGIQMw5XsgZPrIFmLPwwFjN6Fu0c5sGMSAxvGM1R4kxZ2v5tckrXrYZKOxVG6yMCqEKp
pcnQSGB4Z1XTUZ9ETQHCjDUtFV8pRpC1HeIBuGObyQJePBBAIZ7f6nZy2/JMTbIZXdLbp9y5S8n9
jpHyxLSQyaXpSmF5LhMJtm0gK/yMXAzLoNEqd4N1bJigYlpKrHRDjlUwMmRfibADv1RwhNUSQKdn
y8FP8wVPkJIzsl+/z/L/5g5Nc/945PbxtkaBGSRnETmc96WXKMJxP06WLCksnd6MBdZEi5AnTmiZ
+RmIRgfShfcIMxOF17qvW9FPAzxk3Cy+P0WCUWq76YuXEe0JVGtHHb5TSc72wiUWH1taINBaSwGC
eUR/n0b2ms5XNfs6Lqit+TH1oRPE/3beXeQYGdV1ds7WxQNqNKST7Mcy6LjN8SEUk8w7di1JlITQ
tHupKz1gO/cbhZANdP346sgRYqCivnhbhhzmp6LF07sIRu71cE0hEWIl+MKlT7TaJOd9aGcquE8c
p/INnqSZmzQSDK02G89XR8ARoauxjCw/JkeJm3QkBiJM18A1EPsjDRY0Mh65ykqwAkgkrZeb7O5n
iYxKY+LjUdaztzBjOyM5CC7QRt4SI6B4WHI55t8+lxNelTTinsNZ81v3i34nZ223p5aJ7mwFzfaB
anAN+hMrfBnS5DAzFxrf1cHXt+72wECZBYubcA38tvrRQ333Za64vdsXJfcMhadUYc05pTJUrn9m
wo+TNpCNMAygNmM+mLoVxRf1L5GS2eUNbF2Dh3G7rjoc8tTd16jMbAqGms4D9AFU90YAfVovIgRP
1m1pdLb1V5i35B4upraeBxDJvG8HvLkdhFGjf7mUwAAlOSl8ya6cJjm85PtvMkKwf8wc7R50SKaY
S8ta8xlWkdUafKB/Ts54cj+lNKgD5DwjMNQHEveP+YDGviNcJ/LvWtyKdKJdWtg64KVEs6l/uYhY
n3cczuvGJd4NF7DAkjvl6OzsR6qRzg1HmVZlxNCyqD0biViLAvXuBh7fiTWadxBHlslsH2odiKGv
gOicV0KWX+oNkPcUcanSgcCOG3wd3PKepzMtfEhYHZMPiG9yiRW+hpmMsidOEQmgRRRZQG4WaGM0
F0LnH0t7OFvJohpmodIrhVxeUL7j1J+5DF/VHToy9Zsnwl6JamO4+GEHYr7UT6Tkiq+1Sdd70fez
iXf/6fQtQaR9u51BEWkcjD87rl0/v5XOOBayn/Fe6gPsy7s9var2RMUQX3joxNkmr2oHHKO46080
Tih1JgFZsAxmurKojxDJjg97gLZSGU3lPUy2LCcRYdBO1Z3K1Y0O3xBhX5mNj7a8CXpkN+JtBKYl
XimvnWPk+nCuq5Wa3HiMuYDtOU/nf+osIo1boJO8VdFweGKsOvA9At/M5RplaPVwWgv2ybT20h3X
dXB+zSDyTihuTSr5NNao+ThbZSLmYROjnOZ6dvNb56E7dB5GecTXpneGWwz/acnL+uZ/szM8jOW3
O7JB5B+85+TrVxv8Z82D20u/lGpgY7OKGbenGjG4UVDXF2fAlksdALYr3ILXmbsrSC/IWu99u+Fh
AjMNsdPJRJ+OThnrs8c6jDKtUcHslSODheo012aoy2IP8s6cNd+SUMxaf+Q9bKZOJBSMO5bcdM4k
KTdmg3/0wCk0M5MYbWo7MkA5DCjarlmx9fKSefD2a0WcUQTYDM4sIzy1M+k1ldu0BNAPv/+Mvjdt
4wLs7e9vj4cMKRWf/QcSSvvBQCDkDGjAYxfoX+FyRcA96ki10d1PsZ+uqxoCBeeGpBe1+r3w8Fls
xU6QWmXZTx1XBm4wTUy6b/ZvKuQ8D6rdI20xiZs22l98IHglpk69UTuu62XsjA1lgVd1a6CePO+O
wz/cMJSuLnAtHpQ29ofndGcg/gXiV9IPaHyvvKdNjdhBeLIlcA6DRvkpVlKpJoBATwNAQ1UIVGyk
JrfAHg9ubdCbgxywb278ka+Asx2wtJboBG3MqdBrohc3Sq3B9uLECn6Vk8MQvwbzpgL2fpX/jZde
U7WKV7D/lBfRJFZj5yRmGGRJ68gSGV9QhnNWECfRutsVqltzCZdkCbohColnjA5hDFF3jT8lb3pv
r8C/C7m2PcFUWyBjWFqNyYVAF1d9xmgq/G+JOEVZ4UX2KfkFSRiQ0NwPGVkPuE65UU9eTmaWQNYp
UJCyDRWcXIUHQNn2Tjpa629Nc0U8jWiX3VmT9dXIPg4VlOTWnHOVoOPiQTSOEmzaBSNpkpJgoJ/u
YajInmSIRb/F0OnjDePpEuBLR+K+NiEJW3JzhrGC0GUKmGqbEjJVE+uCJAfP1rPp7HlK81P9vHiW
mirt721Zvz1vBc/aJwEKaUFEFgqxRi28SCb36YKFZ6uaqLlzY0+U3Gz9cCXKflOUQOrDS+EH9Thu
4mSAXcywx/8GgZ88hlQcJh3Y5kYopWCwPWwfVt3Fi0hRzKjlQLU8/P2uCTCmMGABZcpgKnZQSKMs
+yAJfCuBdb9j5NRvSK/WUJLa75p54Wv8yGBOgboRNu27BuX3aLhWktzdKAfc+WI1A/fZBLOe/+qL
NyQnSv6ScFbJ281p2eIRrP8W7fLDGVVPJ2ZYhhpY/QaY0c1SpXgK6QYyjFD7ZLG+GoYSdX+7aZfz
QjvCrg6+pZtqWcYRdlAeWTKEm5UzIUoCYk6p1X0J5aCSabbVr/G/OGQzArsbKLmU3hlWa1T9lB8V
YNoMrWJeXTCrrX5S2vEXXlKGXkIgMIOqH+OsZSB/IAYmbG56D8qPSMlT1AoN/0C/JREm8OxSaNIw
GDwG00vv80X7ajuBt1nrRlr6+DvTOvxGxxrlgo1ZHO7Ow5UBt8eWLbR4XfcmV4QsSP96oV7PXOlA
m7DBnZDYPtpV52oxITRmPgsDLtlwy4M9LVmELhTsZ4lgPuXk9PwKCmaTZsLWjPbO0J5MpEg+XkaX
gutFfbmOXafbPfqRByMH9TCfMFOXDTr80DNWn2WeXFDM47Psk71HAbvbUj1+7ES0m0FCpnF72NPK
1NxLKcsGdqpSpQGzlvhoLSU4tnRwrA//dC0+0Bq+mk4DkDnRcLZNkvE2WMt1401A3jrJeQyZMb1A
kOPREMCm4GswUTNllK9V/GjEUYXZHgadj8OPoPigFCTOyi5pV3SkbsqGD5gwIhDiHLr7dLvGCDRn
P7LitbV8LYyEbo668O3VUdNOZuqoRgbEkVi1y3fw/FdNJoGwoT/pblnE8cSHdK+KMFLS6MosTiKW
qHrapaRDsr/vp77xJ70kPycvBvE9rGEpJKAgfrzUbze4bQPlrjwX6GCG9EBnptYFVmQE2LtEuKpW
ryEFxU5Z2YXO9y1e4eOC298y6lPgOr0NZCI0Ztb0ZN5a74O9D96Et2Jcow1KumgfLrmrC9yl2pis
Apz9Vwa9WkVULvokm2WELJt/5Jj8IqflwsHh7tgsWZDRMc1u5SVZFDM+V630XNTZQXNNwq14QNzd
Nwdwcrtbxu9kG/BilTRq/rK1wlvJRTonxKSNC3HkSc0+DZGKch+9uqDkvMMOQuxXxGajp8TdTinH
+rW02ALOpHD5SvwkGMmNRHasrVWSn1xSehW+qY1kADTLMnVu1I/SRy6t4jMG3T88880GUIjJrtaB
iO9FGrm2zMhVXHYnGr1e1vTmrGYGsb0wyOjCJPvJV4k9e+uNofxTgB9bdhxOYe2u4s2rA/W2tbPk
sXvI3e/kTHEfyZBlmcrPKQLWrZ6PaguSi5f3cSY0k+jwIJe8qRYYuAu4Aah9jB0EcvQwtkM/VNAM
pVZof7eF3WSYNU8/1leef5tRNsp2+65kdbfve01A7XH+lGX8J7cf8qBmAMLifb5HFjvfPfgBqTve
8pC/Eq9xUsZ7e+NMbUER6pQWBENazUrH62qBj4CGIpSX3f2IoCmZvoGWYylxnQe/OANq3sZyDo2b
qxBDh/Wk86h1lS1aYMHthjkxY5pPrqi81l5QRZiplwjY79udtkoduO7lPFpKUf9pk8dkjHJpdXTg
ZRx8CDyfARHHUkktKf29J8KtjxoVq4RbFaW5Mm2amyuf8ttNQneaPNwVBpv1QbHVwYLgklDVqlYm
7/pceWhmQMZ+3IY0sCo7i3oiDbRW3wU3BJZNxhhL7q9F3Win19ugwA8Y75glCXWG2Dz3eBfvtiXw
lhdREcPbI83C5aSQ0mZ3IN4xuxfpz9TNzV1NElI2u95EItxOllPUhdTxJuCA8CZCVJizTQDp1mp0
99kCoAzeNvbYzt/jIsKUX9T25T9LuR55spM1WN8KqBAKsWFcsYB9QG5NxWKmUBWw54ogZcZ2wnrA
3IGUGDBgALBrnE8q/7P0FsJt2bkPRxmPUOrbO5Bwk+wM2nVXDT2kzTiezIzKr8mc9SOEPS9vSh3s
z2QVjcE0BJFY3HHkEX09/ymmonAPfCAQ2IiLLB8wKjK1gvHjRU0eB2yb8D7XdseCIHIoyMekY58F
DoNmZm1Fd5NIgAjIb6B2ci/8IriIi84cILGSg9s60ovtTm7Fi5Kbkw9HLT83Z8BNOmp5rwcSSSBW
aiDmzfoOPsBhp+tbeMEmpP09IGvUaeH2wA/Dk63a16YHfgw0EROeoFoVc7Y2joNJHGhHuz92OJGb
6PAUxK4UQ++GcMPe3+dY2p7k8y6IeCu08HAZ1aZHXs/hZ91mbmISZ5kGvejupo+UxUtxi56jJqsD
z9Xt41WRVFK07kEaz/sSwP1pqWVCn9javAM5xB/+3FUGQ8/+Y0i3ebQNoSbsCFnPTcxy8AKA7ZDG
DdlLhEE2sx1fG8lHxl9geWTTrWM9weKGf9CWP1gh8eIo/U7JiB6n4d560TXGLNt+6st5VltpKpu5
Qe5eq/SY6E62S4sVP07d0eoTr02CiqoVTeV/2gIf8HeqXd13LPV0YnCItwott1vSzHPJSYJ+O+ZR
jWSJyLb8PuW2Bs4FPAx3j6XB74vj3JkEM7LcVTzeq7FpHXsddADUJ8r3HGooormIZs5MUgZXpebt
3E2pEdJDf6uCeuSZnwBFA99zqcYvKoHViTmVSoavgPeCFoPXQ/x7snPFVRWbudsvIpYwUORrBm1I
H1sjM+nLxk4OKaLpfKCpsTVB+LzZoGZ8QFFauqQouO+SLRiTwyNnZYmbPTzMKm0VGLXSgUsC7Erd
ceRQxDo2L8ENfheCrjaioR0X2NXHZlyYSF7j+h40CfdTwNrGEfCijMIDJLF47X4GP0vwyvPx6foP
yPjcwgfZmzmZ97gS0X2qMATDeUcD9LxIaNZpSBhJf4a/N1iUzSbV844aHcpgj52RVRgcm4vUX6PQ
LUVf7F+UdqhS9gu5/dtp9gGXYW+mx0j60B+Vv1dInll6XvLuiFmC+MnBYEjKiObQgidjf+PZ3qMe
mQXwMp7U6QmBnIvXXDsHJUM+lGsHQywk46sD5F0BgVcwENq8syN4KCrj8Hk24Jj4NaAL5pPo9bnJ
m92duT0mZNvDlg4KPJYEQE8xCDn+AHPzwDi6L2UtjMDFFk9deK96PH1SxfavnnFKgAAx+lQ+Ijsd
J47eE9rslDcM1V5GLBNE12HhLgPkUkTV+5EDBmKRqRusQmToPNKd8665V99t+i+sJlwpHoV1nMEd
R+m5eBbaeHEwWS/tTGV62sGDGDLLTSO6h+23ILqWCE3zDNExoQg8tCARxC0X0uuX/+cXZ6mnlte+
d+WDOtlIvxiF5Uf80oLwQHFHpDbE2YXCzE3K1H6QoZcC03nH6u21pdYpik7g+SRdUKEtNy5F0FyT
nETjgg6p9r/BNHRgEY4iGZaTfSfI758aAXVktuknbLYeb9fpVJ87MFvpK+eEV/4nZeSV3Bi+RF9i
Mdm+rfCZ7NQVKQQLiKCHKGDSnZmj8NUCeKuOZ5hnGMnm+fwsyeKqlS5oiIFNbWxSEWJkjjeSFEsS
5eFnFDb5i2zZWxGGc1yNHwXH35RRoNy7LaMzAvy6gTqUNv1xeL9ao+gXn+Sr5uWQKy05Die2p3km
gJ2s5phjSmEf4jyXLRl7CX/D2iQsQtxbBRpmNrhBI1S2slyxj7LXQE4PDHF/X2zNcIVyafzwPfy1
vbMKF6LUdXlzItpn/xt/IJ+mmitFia5hig+D5AcUKbZ9Ey1Pwwm1/c6WhmWeuniAyKndNLpauJBa
lzzqASrD+joN0xbQEpp1yGG4eGz8prdt2PLBH3V2BU2RAtMc1uSJ1dpX5MIBJL2Z4592heR0stw3
tz1vtlt7aEqfdwJ+8EjF2C8O8DQJ2IMtf8B5S4s3Cv5cjSjKGY2B/+ixTHdzMc1CPg9vIMfiCZVI
5gVCreDQRKJk7jzgiBfUp85oEVNDZXn9OMquydhdarYYYganD4AN/kfXOc3jCY15qehg47Nqaqiu
KSii7sk0dR9i2gJYwpSf1B2vtm04eR7Cx3dlSVN7OXrVEJyZfc4da0srY1XQSSKeF4LCCGIwy7hE
Zau+tcZDjCDDs56QTv6H8iWXpUwEGKg07u4H32PszYcBR5cfY3izFDUIoX3s8NdqQbXEZz6dt4lx
Za1oo4dqZBRV6yAiLKBXDF43WL9vE8U1wBg9A054y2OWgonzUH3YL0zI0QZY5fh8yM9ks1NUTl6t
GR1jkJMPpte5Sopgx3P8wLMlk5HI4fYnwDZaYwFrxMNYCylQypQM4MgH8ztwekVoBMfY+is8Xrsl
GXf5idZwDBaEYcwf9tc9t7/GTiqWU9E/ynDFVqN3tQl4QJ9NwudO/jH3SlshdMwVU7PwFSPUtlil
NWp/i2AI2pmdvuJwaqhqmE2FJMzcrybBcKS7rEZnqZuDqP7LDhDMZ86fvA580pNHROpbZVHU1f56
v/s7E5OZ4QdnosiTh3zlUqg2bM0scujBoKmp82nQ5jl/BVbBWbAcLQvR38sP8eZPIGQv9XCRtIkV
h0KjqlyDSRYP0bu0B4wzfEdMUSLel4AejKzYV3IdTi2uDlkxL8EDmo36ViliJ4wqAFqBuyPDbXbk
pJnr9T2Ui2ORJrs4GYmgsUTprX8oPKqwYnr6l6k5EBZI9K/TwF/SHRFjbYK/VVg8x/fz3acA32YR
PjIm8h458jeIazjejkjxpsh7E81qsHCx7x+qfCYoQ4apStf8i9tQdnVhAv6+0V+ApDj4cBh0/S74
81AELK+3G/PZAvqGGZxLU25RPEoGiMlFD4/qxTcYy5A9tHn8WOuM/OBY1oatNO1oMk5L1iqFRTk1
vA+WWv+SvtSA9JiM8++WXvj9/skDon/jVBDGRDPuA8zGjd9cu4AQdz5YbDgTQ0dYOio3owYMkG0u
3XkRDsFjePQMgPhdraQwtlfzg4VUwWKSirfeCIXQnpj7uhvxuNkY8hxddsxoz4Z5v4vP3PQ9pGB5
n51T31bbcARvkBaMPCp1Zp+dg+e0yraC+1Uh/Wl9zwoY1YErYh1WBHIUaev7aEexvRrCkNCV6BQT
yJp9tRlThhmyMv+kNu2oEfNDgEEQ93nFn7UdMqg+LRhKSqTr4QgLN+rLPjhKDcQgbh/4e0nHTRsM
vDBEcxDCtPrgNIYZ6bLN14lwJsGwlI5jBOJ0H0GXXeepjayHrMd9LfqsKrwmg2CJY37qlEKO11hN
limdsp5xdM/MMVAFv4hk41QijrO407HE1Tm73CB/29zaXXoeCn1eYSibmC8QdM1FyNrRK7VUirC4
rmTdhqB0jYhdvqZeekGFPwvcb9RVJf/mAfxwgi0OVy6Ya0yUDq9ShFxg+izOngRHicVGNkL75gtJ
tTv0McRIb0HSJ5iCF4ZtzPSLO6/Vpng3HzjDSmEj5elqygIFucPaKDhxuNsLuu94XYboY7C3nTzp
XvfgPHjuIu9vtlN/S9XHFbeXBj4t8+/1LGXypjhuC/n+IHCVbTY8igq44p0EsIzY1i7Osy4i0h1a
IWPakBQU0oxekaOtTrAYpngZOBpmquYD3YlnVm5mldG4y60CnzqACBq0KjniNkdRt/zsEKAib2Ix
3B4CpZkuwX9JKk576yPubFbP3aK1YJkx834KFajcrrLWR4zh/J2oHkry38DcVFWs913OJqpoTsi4
iszdlmSdIDXHSkLqLQOoiAgyUorK9y8qkIzZ+CpsHA+Ye+k3fy9A2neAYSyXN4Os+Zu81JhirpeH
QWQrL80tJvUcokWXuX3AusORwJvN6ortRevEvoMeu1lnssQixKpSDEiwfRzXkHIbs6no+4+0fqpG
Iw9AAdXolSwBSnNAbOXnCHRsvtG8IBXuAyg4lA7sRhZzYJULV3bajojI6m4ZjZA/pQmCvuYj/w15
pisB8G7SATZ9FExai4BBgCUEbFjvGjJ7MFa97x1rmfPEYkfZtfUUS9h6tsKIpaLvlzxYs86PiKAD
3HBB0O+5QymfRmtVAM7A0PtcashEfqlq3SYdXPEgaucDADOzow9NyWuFcvQkgH3wkKpgfSkHjxrt
57zdFympX6JXY5UN+++fggCa1+eAnjvmU68Uc+RckBrILh4I59dJ7/ENZQZLSpxWvnvKzdlXmqMq
G+tlI+hkSUiwar+5lSuxpl8ktllq7yTTiRW55m1VvvdL5uygKAgCXN5NABLiwegFLL68U/SF25nQ
bR7Fhfdx4JgV6dusR9OBwmjg9bw4ymTwcM4qQ2mu4vrYpuXtHl30CNcx2TVGfkco1q9iYY//cHSC
QQlW2vTpyf+f42tEDcT+/xz8LZzs1odkP9wqe4U1z0J2WbGvhprBqXNj1C2rncBZpdWheqYapB4c
H4Sn1TfU+xq/agH++zdXAuUt2LRePOklt+LipzB+EevA4z2oIHl447fjnha+ENgRHuWykguQX9wd
vLXhZyu25VQyuoROjV8ynOf9w9b4ogib+Hr2aIppL+TdCnCifRvc6uzRz+0v81Z0g7PNujkJ9y6X
wcYrpNI0NBNKnnmtbGsm4BlE0J8NbcLTduqRcjGLsJY2MyHC+9nYUWgyFTGULugzwgvw4CPhhykc
5U6lSMpjDI8IOKYExlIqMoXVjWwkQNyoWkn64jm4eKpFXt636WwVqNUwuHoutc9Ym0UoIXGFsCCy
KNXHB37tSgZ8bKANRCmO9LUp5CgRiZdNOtuflxsjBPp9e2I23rdEbN/aieLoqW+1fS7rOzoI8bdg
/NMGnnPK7Cgn67A9UcfLpZLidhsp7IhrIng9F2Am7sDx3s8b8p4eltfz+ha0dpJuSCoi3vdmobYQ
ju8hFTzlXR6Sv0eNORNuxlGvMz4Ag1rXTo+AhGbaclyBHw3qC58NYRk3WUeZj3T+zCUeAkWMMqDB
zcrbTvSAlK0/XV3RyQVrhuyQzcRY2gaHDBMTV6bctWK0rcuWbF/UWWpBibGtirG1DET3heYr1pqU
ZMtAt5iye5644Gk2M4dVoW5WscLQhFZTt6v5XSSVjG0x4wDWqWqYZ+2EZhqTk6FbT5hXgsrcFCfc
DQXabGQoVzUsk2laT6lEhfy96U5fEFzIoAuqh16OmgzX72ErNvUoGriBeA0J1gYNwdoKl4h4WluH
OABeaErBeho5TVwTN2H1rqb0oBhNBXL4b8fyF4szuEejFew5K2NSHmJwOGjeo32mXmK0MVwPa35P
NF7uwJyE3iJjPHfmq7wzYs8Ib/us7mM5y2BMxHjOPJb4bKCLCbwM3FCfEz8ACqwj+522Yq9iM2yi
H3NqYeeTYes+XnvT/QC5bf9/8FusxkXzrVWo7cSWet+wbHDp4pwXP9o+TiaG0RUxgjpkc8Su4qLX
5U2Ie5wKyoD+0lalMkUV0ZWGTMSc25RH/bLOxhS2/t58Z4K3SiEkpDmK7fAzi/kcn244XtBsBB5T
JUXsxX5BrTvvAvxWd1ui00l+zfEaKOVuWRfsOxV3ha9Upd+rdAeOHEO1cNIkgA+yV4DYuuPb7HHC
3r0z4VDTvZJZVlhI5JT8dDakTiOetbA7uXsaWMow8JWVXhBlfIEzqRzHk6blVV6mxTR5EokaPcCY
oyAMwblakq77dOld793aqROw+hexFQ95qPYRyzfJpIIkZBQxt8i4ARweD4dkd8D5YLWoTCv5LIde
vDo7Uzd2uSq/if67gSgEcA1dzJySFXUULCW44UYk7Vv35ynXLNScxCq4PqjkvUq2es4n6znsSPrJ
zR3wUBXA51IdrKCGGHQf+IEN0mdNQOQTgWctydS4buk4+O2x/pTlEJdB9FA7G656M7+SK4KZOr3b
0SXvmYId9V3MypOppn7kujRomIBeY02f4NeDS1LdpXC63OQIr2jxnXJJzANCvyPG57NS7iYKXJ8N
0KuSXXXBxeign1bkA8zCNlpbVOwzmTv6ngkTD6QKcm/0PJup1HT8LTiXK5gEECUshYDhv98GEYGh
Wav9qKGdx34xulnxGb96o4cKoO860IjjS35XMZv+ce29bAEaMPb8WPRkrFetrZHHPanMdMfZNmZ1
qIBD4qHNiyqH8Q4mR56NLtoqJFuPn6WxqF3x6kv8hng+RdtmavC2ms2Ohi4OuNqSbfZzErZQKWIq
f2e0nP0GiS+tKOgEvdOjKpD8orDxjoifblqUnxg7ztH4DmeWQuFMErvO+lAhLTeARNyS2/b7uT/C
b7utup/V5qadT80dj6NJ1Z/0c4xFmtDW6CMOPxCDc5R+C6yaT8ouXWhcLQDKIqqsesnf1E+qsVHE
5uQ3P8X3ceFFkzg33zQZIqFu2GEiCxLIm5v1ZlrypTwVyHULLvgv2LK8l/lSbzGX16yJokfXHMgM
S5ySxeo8wPHaxiq28UseIkBE5ZIy22ZH6ukJvwcR6Dq4+3/+LwfFKWQLjkSe8ExOfzfTVlbzTj9e
PDM2sKtciownGdnzifEj4bXc7ztBuMtTcBbCcmxu1ioSfQy1m/9aVGRKMRVqZPyB56v+PDHlzbtk
HACWJP17Sv9QnEak4/Ari8vowovyW8hHC6LPSXhV/FUqC4HmnttV36Cv6Bm5utM53TlhRQqxHClJ
zNc3jSSpb5lJnPkwFcBpvLXucubVziJPTO/oYKA1lIDlpcRglNhOYGgkNKFIqwbmABEgK/FLvd5Q
BoK5J9EfagGbMw1QGTtggmP46ZWr+nTU+5bk22H9j4ipdUpSQOpPcMSxvjO3/BiNRXb76kgZ17vC
KE5ZYOSDpcjpP3o/+YWFSYZq6JZTBUJUEpRUSEQ6iDZDt0cT4JgrcPHkbEeTdsPLghw2j0zqgdgD
gZJVPWPF3QWdY0Q3VFFTm7+8v/IBVkkBfLpwT6fyCEKqOV0bZ3iMDgkktdB7cC9Ww/fE9xE/WfDc
8mc92rfUqZ7HBDMLRxeMeRKW6d8CNUPytC3rmLlfQx/XVHd+nL/zvvQ8vRNQyotBRkYi0mPnVXMO
C9rSu+YUDx/pUBmMd1BMBauELCIRyKlNL/laLU+uwzyjWueYsY5IAk9Kl/3dvnMcLaRJxmlwSGBM
Qt3a2DYREjFfgJXhdEXswNQzxNn3s6xP0Yrg1qgM/KRrnk/V8csTVezQi3dLWu1o9EJ+xOLPgjmT
ZVv7Pkz8UgQ/Vs0Qg9feQHnHb4moBVeQL32WRwlX2/VUPlBTtLrXG4VILT0cAkQBt81AxPxTCA+w
5ADzhjyHK2/gmR5RSbOoH91RM0H/ewHQz51Iciua4tEwYOrjZJHBunnUk4svhIy5t2dg8bFSzzWt
qu/YKUhwLCFP2vya27R8FcPgfvgrD2JlMPmfJhYmB8SzQX4n4MsG6IaLkSL/Ltk5z+SBMt+C+XnP
Q5N15v5k38weRs6fjv3T+5UFM4JCipmMDLMCCxu3PdJbhAC0UbD5mCKkgMaM/rSQKo6X23IGrkls
FkEr+w8AnssOSW3Cxg8budXkkRvQVzZT5nyMcRGRN35gRg8zlqF1ZXQz+fx/zsCnhFPtxCE9Ch3E
5CEc8MzlezoHKc9rK5Gpkj86Hy/SFXLVYP8Qk0uVmLJYMqrgE8+qXAK9LhNSGxoLPOYK93PsFuLq
h+B9T+m+T6bUums/MGINUlZESmL0S7kQ5qUKn//0DuPQvJSqDgQPjgiXWuzzIw4u/n9MVkVIi4kW
Z1+Q938LxCD6kNwjoIAEqQKjpu/1KlnO0oipIH18CLXDe1YnNs1e8kJ9PI+VcvksNPSpRlfMlYzz
F6Wdf9exLmSO6A2Rxp91mMUbKdTyrIP5G92W5mEvfOpSUwthBTb41UrS05aHca3AYxRmZJ6SmfQd
vQwiMraeRLl2X+mVOW+++6uSWodO9tegO9oDhXboFkiSt+kTF4Etkfn0AXLVmFxbJOKuE8MfB5c7
XXGRGrYqmdmztYm+HcNjXvh8gZmDKSPz1B+1Y6qEBcv/5Y9onu7exEh8rETB3miW9Kw3KSNF7cAr
AcJ5zR4TZW4ZOZjxEY2gb+LCIab5M3KZ17GDjrs2PCY9caizv1CN3JCrmK/Us1gVCadxy8zovsrW
F9vG4w/R99LLoRcoHmUdMx2f5AhiFJQ7TRJoyvTuJKFfO5h9AKcRIjb2PuhdFPXgJidjg/XOirCE
mp3Gj1bduc+oHnV0cShThJeBqerUydnJyv8vRBBACpDlzJUZTtIW7HfKqfbeNRPOfzDHNa0yt5Mt
6KXRi4QXNwQvO0KmtTZHA/YdM68s9OdjSBunuUIv/GpiwujN2ohx4jQoLTq4+R+RGRv2JnlenPei
frwUFE66e3/Qbm5FQvI00c53X4H9dY+ORBPr50w8x9z9GHeUp2njEsrZEIeCyPBF4RC4L6qtZRDn
QaIYYBm9Ks8zLsoqCiB+u9t2LC5knRFRjPKV2ikl/QLxXwqtr3Drbee3hjDsvCTgUJFVcDj2xyP5
ekq9phAPzSNsh9RJo+OCppNU1ONcM7U5isgbtVLOIaSzyn4gTu34c05l3JqEbqAsqVUuK0cnVgfy
bzp+zQAfNV+Y8M7R6X+PA+mWjpZsv7zDppPREP+AbjkXOgJ7JWO4myT0OlJyd/NW4NX0srbtpZ8d
8a1LnzTD41kj9cKE8n9j+97B34f+jYzp7gQ4ZHKI0qHIs2E4q2LbbXUPSIGyQub4KGj3263izhEg
x+TqUKaPc6gG8/sKyZiBsF0ImE/GlYrmGn+xqS6gfnxlHU8zfg/VsAF7IpoWSOaJ53wCk0I9h6bm
le+39RgNd2BRMdXSixleHIDdNo8LfWLCRld6CaWN0OB1J5xmQr3nlggQJEX2RT/XMjmRRT7TqyVc
uKsulGxnRZ/s0FmLtQ1WpIKItCEi2p20UDgWXFvhQCgJs5AHsfFimtbEEQLs10BRqKrL78cjxt9R
Ui9Ht8RR+HdJ1s1s4aHqdhaYxOpYHUZxvPjuU6n3hDNHLj+J75Li62Sm89ZF4sgwUSdp2Ch1sXRB
vYuNLrZnrn0ynGDPmVDtWvrSIg9lbAd+8QQpSNxXiGcMaR9+kvV1M/2CaQsBfpBrAVa1DkpU7K6b
hqPsotTS1fdYqEbN1fH3uOkON6eGuvJWrRX0nKPr1HqsAN+eM7wtMoVVms57/kRWVVwsGfAQ16CG
j/dPaZQ0Nge8Lp6xesHV4/Jyqxath6kJvldJTI4l4ZvAW90X26cAxtxEjqg8k9PiZwVuhLkM/mmz
UmQAG8HVunWF5KDAqNNDgRfo0APp7Que1QJCl7L/NJQz5P8PYR/+TqGdT6oqDD7jEsV9v9N0wqCI
AF9s9yhW0nb3O3dpVi6czLQokN+8Gf7VNxkltUbaqTsTz4UsGuQ1PQJp00l19sITCNz0UsgxzAqI
SAAhSSdBvLxtmCcPW92FmEBcs/3IXBa+e+FtzNRwWCaiXpaMiADwzHe9YrTw3pvjMCBljeuvKGpO
RnLGQ1bvH37cAQ5wgF5GmKSGr6Mc6Bs2nwJv78DR/aupFbMjPNDg8710iaVu/LZvUf8PDnQxsN7F
04sCHCEcFKJEA4+y5oNQbnQIuly2JKou421rYdUXQocGqE8qp1UtDvP/Kqwe9OEU5h+VDV3xOAjW
NzCVbkx2FtDg4j80wsKlhOyH5cDsCXboU5Z5JgMBmbAKYWbnpLN8fc0nersTrVyKRYKpM8zWFzQf
WaTTGF8kqrqPCEM8lGqFyd0fdI9qK/XXFIOifqBUIkBHiMKU4k6JTUxBZxTdgZHoaCmGwLO9KJ3p
fqFL3ECehK+C67Ix+XwTWqhnRpA1zIShLjnRaaMXFD47zKjzDcGMUYAayGAIKzIcHVbu9G+/NrRd
9k8yDivB4TFZLmtJDLD+Ri2Xmkz7T/dz8PHRmAM6ZhTpnYQ4lUBvolmBdHoN4Dx1mhN5iFtY9NmI
MRfelL2ym6KfUZQ9AXy/EqUNdjp63c8SKVo6m1aGLpIm41TiioW3zJPXrUYonEUu21J9ikvtVEWY
7IH4vUv2ZR3OnD6ev2YIRO/3+uO0XuF77+bxY64axoGbidRzYS1lB+YbLBvKI7cvLZpeIHhslYcC
MpK6OzPBOhMgWB1VXdzIeZnswm3pY0JXElgwFvaj1mGLUu71C/zz4SNinP7cZZRhdacJx9lWCYYd
PSh9Tui/MI0MhmVBkhQAb1V1AnXRXz5k/3pE8fur/5drWVFR4IQ61afME0BwcNBqE93uHW3uZVNe
fFncJSj8q9KdNrpwJXZiiJh3FP7JXrMOyTRst/MyrFYuqzmPBFVBAEAgsvIuIffeeLsXXY20FCRj
9NS9yPOh/mhhBm+RNGkW38/wHlIFW3LG2sDBfHxbUJ+drjYnQZxtkk7PSBvm1/PtZFSvtrBCMQYZ
v1/HlsWogZJcZn2HAwvDigw2YDaWv8Tz700qOgP4D2L23K4FsDk6L9KAhJRW+0PQ4lf3kGDobtsn
3AMjaDN5Ntp0moZ2pbZPPJjAjo5/DGyXuO9Xcf/ccrDNcN3xVNrggV9J8TtxxPjiRSD9xhB8pUS4
qwscBiTY9EifXFp/gxF8N0Mzg7wV3iqLs2ZvX0LtjdT5tR4/omRJEClIsNf5iaSr5QsEqWqcNesx
KFa1CDQuNMNL+Xs/boIzrBPjV5t/unxvgpBcGj4fEO1gX1Ti5etEqm+khaKWxPBZvxFRBiI4Krzl
v7dn/KowpB0Wrksd0XUkT3BsEiiwrWQDlWfWH8y7czFDKN/ly+6+uKgqu+a0I6Rr0XZHd1M6Sc1N
87a98zBBLVKziyWUQw6H1BpCOJg90IsD7er5Ic0WoVZZXehO3TtlOHWyBFGGZF7WuVFtxoJ/O59q
CBNym58o7YpyGxJxATUPxEAMw3r0OrfKtHelY9bl1LtFn+WQDIAUcp0sIB877L1lU1jYmuCbSazj
r8Zkb6rX/sXuYlVgNMXfMt+5Fsz0bphxVswDAAyDczcExvM9BIRjeD9Lhd3mhBVr1I0/s6rk97q3
ZWHjPEkQWzUnBYx7QAGICQzM/+owd2omHa1E/Rrws5YM+iDZzq7gd8Pzq9LSGE5JzA3Qrg+ptLgw
XEy1vSfuvSrSBL/VB0DSlCwjVT1OtMy8l2COFB/CHSPk4ALvAK3SzLL3GHYXx1JR+xZhzDp9MSL3
XbX6i9iRcoJaa3LXX1ZIxZtm2ER2mQQYCFmf/4CRd75/oXSHxyUKpC1uGq6TCeZWi2oM06FJPk5+
Ll9NTpZe6lCVCRlkCYETbFfcQbqkaZ4Irh4wr8aXmNAUKYoEaHQGALVQc4y3sCGARgRBqOOj1J1U
cBJgKGMj9lkdkKKbYYcU3rFSseM1F6Rrj9h1y534rqt2c4qCvk7qzICOMxerH1EPpIDOYElTfjR6
IED+ssuWRXHP5E+fLup5RSAJe8PsJ0Odpzlza3cLbC9HlC2glrFfMBF5O3cfZOKwFmTL/F3BY/R9
NJhQ/7B9vAy/jbocydU4TNGJqqhk3z1oXLO3CZGCO5A/kys7Vn42oCemW29f1UC00mm98hC6XBtH
XEbAKOT9Q2KAGkpcdeqba3L7SW2mw4wUrhvlWAkBt2NCtF0vfmS/m1K5oBWZMWwMaG7yocwD8sAo
hy2zREhFOhQuZ04paeEmI/YZT1oT8GtKq588ixXGPcEAiZHDtHWeQofj4oaAqzZ4auPSghB4pjOO
cw+kVNG1oRyNyf5Xl1DeWZPUklLj4pwxq3Hz9gCzdahVPJhyP2VFgdkoEw0FnwLudhRPRLjgALly
f1IO6+gycJesSGYn9dAlQxXdbwNw0pAXip9GxblSyFZhvghethkLKbUPg+xo844KThCKncb2+myy
MYKFKAhDbTUVQQ/MGOIPDwODol2GqpujRq+63w72PVpiNKdxkz1QbjIxoe5fR4zEVWCq2TodRbNY
D9/MmibQTm7E2j1Z+bFxRmG1+SYr+6zBH1VMDV8FOTFAv8lVkWqEKbfxqnUcZWGH2qgUtzhaBQxE
p1QEtUj5mXC1rOHD957hka9oRunnKw1NptbBJLKEvmPBxGGL7+CGopnwxjkfmeebfbHWI3xIT1js
4KT0FCGn3V/WpJyjv/gzWN/PT4FcP48q+B4/s5IR1kzSeqRJfc/CAqoRA4FxxuoAFDvrTutH/i56
Atfy1O8ffyCrIMaMeB2SyPewjxT/ruM8qWMslxqds6AS6Y1zDO1z0mdWc50Vyb5PkPxy9UHIMa0u
M+I02rbDxnhgJf5k9ObjxcoZYwonJ9V89nxZPdj7e3WtPnqOT/+L8+vUB+jgtCkaGNybycWVYFoU
JwR3xxnToQ81zNFmU3e3HOJFhVy26BYi1/wSmxLV5oGNY46L65gPtD7JLAbyjdqT7v22jntJBwHJ
WhnRcSRJ6YtDXcEVsbRbLLqYhx0U2j6pn0aY0KhO/Fpf9Cz117gblAX9M4zXkx44Lc5KO0V2GJz5
N9MWWFXP0UJbY94Luxywrns47mxPC8RNMHCVnkgxTMTVLNf/hQIbH6/MmVY3ESfmqvCoCMpQ2fMs
BlBt2VonE1+ET+9NUBmcPvf2vFr79AAo5G8F7hKBYD7DBiVRa1KPCWykdm3ZicZ5v17bdB1AV/lq
zu9HxmhrmMmP5rBsbqwLtJ18Zzeb4VOJuJz+bMpaqyri0bDZ3SlVHCuvpalE3AsSbiZ7l7ZlXiP4
iwh+PiGZP6JsbryW2ktWgWhhOsaXFwN0RVKNlt5sNKrH0NaTMOhkSfu6h0JxDNiII/iSvcrWXN64
/4ftyq5PGG8Cye6DYXxQudqYRES7MF/71QAwevOrL+4/kDc8KmQXkmJMPHOICeMdiw/5Yg+MTem1
Yma5JNDPWwV86k4WA5OawA6BRzEOgPrd8X/m1DjsxJ3bCw/uAMDIv+Pje+C88z4+NUwluIdqoIv/
oj43epT+THwm3GZm0KtR8nXWV1qyH1jy6VcU63m7utWbJRxGqdkYhdcko68jfGIoj/oymatn9PkG
jAKsJh8oJN/GyYfmN6RYtM8HJRGPMCw0tbJwua0bt++OHhdAE/55TR8tWufLZ5TZNmXnTsBGdKpo
UNlFXJpF3TFzvzLuV52tzh28C1jrQ797y+RjFTUsKACa93LozFlPq0zZRe1fvPoSH0X35N0NIhth
pP0ZlwxN1nhqHDwF8W64IVuYX7N7qotoFn8izNGFaCRIsrF48yqTaOY25dfYBu5tvhx8xKm8SfD9
p/MNfY8fOMTi1PTBrEFUkMTFx5aIcLkTmn9OzbI2cLt43kPTaqVx7ng/NzVRKAE+qtDY5rjwp8yl
U2+WAYINvO4PLGAQeE0GW6BhHALGuu55VGIFW9EDoXWzJFafYIu21i7T8/sYzwUemVW9Ij3fTQpn
emrs5sNmPSEEkNJSnqGssZ0mecHDjf2DJ4kgIQq7Eso9UvlFx+jm6sOySlg/M+QIQ+zpzl2gCHaq
8RIMXp2KnyzIs9/3So3O216nrmmWFg3cJLBzBdosSXmCrw0Yko5I8W83ezet2wiJKaZq7c2rCpCX
qPnaxPbQ+8xZF+Jrz9PqkDot2ArPqLIokkdOkis9jsiwVMCkn1kB7pXcwNKHtavA3FnLj4sj4Loi
Um6/epF9XQ8Re7x8AL7dcpBr7eFjOvGqWQCgaxMmBOsLxlpFb/KkP6aihOYRZ/WNglX2OZHZlc7T
lCN5POVv9+2tvkZUoOieb/beYm7LO91dfSJkZV/cwPIh74ONUVNWJcXT88apPLZCT3XCoYl/AWMy
NQMOQGoxCIJVEivexFGy8Z03VnBOQq+o1DGMf7XG0PPmGV0zbOma/4xc+JzvUoDNHF7JxZAMBC/z
iipnpmQu1e7xabMdo+WTnHlA22b3Jae7ZztZS3GrSJHyvyichIWNXBx8MSEGHhR6umYjgyNJhHFX
59WWomtYDjsSHvqHWf8DrBSRsrqvwgPp9JcqfpeQSqF5F2Qscc3nkOgchXcgliGKUCP9Sxg0Z4oi
i+Nb45m/6Da9Y+642MJgvcgv7yrhAdHbUF+3LLH+vJ3GaE+ptJisZUnkJ6EPiBIxaqQMFHvjpETy
0K7Zx+DrtyGSKvv51lyj9zPNVyhPEyvmyG2G3PjA8bKrX1xCKi7yM1CUn8PWqhdYLdEKHlzp8IKP
pK+ra7VU+FWZmYaJv8fEdxhafB+zrAYWm+f2s3RTu1eW7AhadeE6RIF9zbsF7piMxlY+pyPbsFYI
iOorGMgbutr0WcN5/WNrRbG67v2f3qHqX+ObbyidTHQlgm5Re0Wv14norAewDGbuR61mcwx89RKK
wWma9PDXk743qydKW0PlRFrhR1BY1nCuUHnmYnWONP1me7sKuP/Oh6Ds7ImavSR12EO3oBNAMk4H
XoOzkv5UFkeTizzqyukoz7yXdtHVikrEt1S/kd142+ifbLVoRpwJxk8/y/mOZoppSy1ZNPYXrokg
nRUqCEby1Zx17KsXy4psLBmlNA082B2HFy9R0DvlAi/ZnBfZrXGYcAMldAe7rumG4piExni7RZXt
ZGBkq+xmQ2exnDU85itrdqUuFo1p1bz7Ga8RbaqPEj0g6Y6JWb/6tvxx0ngIpHvueCyN8n4l8JZq
Z6nV9bW3rcqWNVhxHRr8eBG5g+tUoPMuqb3CPfRJ+swQZqbja/ZD8SmqFCOioBLYydwJPfaNQexj
s0VqQWghQQVoykDDRbQeCkzVQTkT07TO9Yvev1H5I4FRcLUyZMS6+zRUYD448BG5FJw/8WOrbile
QwjoUq6s4y3JtM9FZfKF7A0B2sU0qIdFkRiGGqdnSYMzIlhqttz7LvqGpcWDf179jwuzE30TGAxp
D/fdQC1S8+6is1LE0gGweV4D1sWmVW8+swXLNW3ELcehjkm9qD31kOAILWSOw+RGk8q3yKOnnRsc
Ma74vKdQHL3/C2dRb2G3BLgQC1k4Fkj8XAeCNP73ROQ9Pjqa7awTHa4mS9YULvfgFBJC9fs4o5UQ
ux7j3xp8LzlPgcqIe8EzQ4zbDo5n1KZ9MZbKrmhbTxLT0RT6qBC4MddpvD8RQ8hS/lpbweEeqIYc
5OEuTCjUyL27SVkHOVcaf+lxkQ+OVh5dhGs3rn4+9mUsAyPGIEcZBZOVwcr7hUQVLCby64IF1W6k
nh0BbnCI0yG2MPswym25v58o6glvomuq6my+tr9TSF2q+rjataGhafKSl/QB7xELy+bIovYhWq9g
VPmUWbOZnZX5T0s/GNW7mS2I4qAkDI7oM4pwKaMnlQTGRtsT53AOLCzvv52hFKeawQXGiSxfZA3s
jXtpqjxDlBZi7LdZAvuGu36yXPG7+e9l5JjekqxBgsU/CmwhdDMasxk+oCxr1M+DGAoytVBfv7lV
FhegSGlBfGJ6rjGBFCyNgSDE4LyRTXJGcRV2F1ih+MqYhQXDxIE9dnt9Ij3wg4h7rctMY8Au4+Kb
64xis4fQ1nDjARPXdhSqlidw3wJCNseJXOjC03J7wz2ssBglySGzZYF4tHCsd28VAvUpmYpNKxCR
AJ7i9cXODfMCbz9LbjsCmVv47PvVYjyoeZdfBRNcghIP8undix07BCdn7TuYqy+Q3niU7oSLKiPh
O+8irqbvN5/vrrV07FbvTXodYHuI+JaaX2b9HAXt5UdYYY/lFF/frEeiWd0F+FJf4Arfl9MtZ9JP
UnJXTnCfcAYYy55yinmU66BmDUuCvlHlx5QhqvLwhPQcAz0eK07FSE8L0rYn4fdT3GJ2d73MzaDy
H/rrGjDT6tkWihOeJmulzb8y4Z6fAT27dBfhqRagVqOeFpDCfzbdHJujEjiTfif8DTaORjBYlliz
+U2ZZQ617en0kV0EVRiYh65gmwqW68E7RuW3oGRrl1yN8vfoVSv+cDGbkHpLu+NrQ36F6Bm1q0DM
XGiastigDmWmGZ0DSyYzg2gHW1FnHDChqxIQgkWIj13RYdxbcJWPD/MoEoF6ltL4jPqOmMxNnhD+
IMrOxIkdFLO/d0qyq+p4xe02qOZClJmDEW49tu7AIXdzis4GZOglWiAyeM9xs03Bvr+gh6SorAg/
XWxIJpZOlKtEaja5zM1Jx5oxfhJNEDAp0UU3uI6hsHJ2L5aZ+PiI5msvJithMfdmieJuvhCijT73
p2fyfu5VC7824sfSBVXeyLN+O0ucbEvak3L3HPYs8WM2OHqMJ9r3enE/2tYfQUUb3d+ByoGHWBfg
nTh+4Y+TtIWlmkj6+tno/qwXkKVyRPI9lHI6e6olwtuD3YLRWP9jyk/G+Qm7lVgII735Vdy3sRY/
ZAOfm1dGo6YvjQPOi0Lc+Nhy6wO/AvZ+Gn9U2six3BL62tff8hZUIkm6Hks4GT4QmoQifShTWNFD
ZRryPPNM5+oN5VtHTqmLc7OQOfoL7kHI4Rpj8lfDWoOhF7PKaUTRWyugYtDL0xAeL4pjcx8l6SiC
00I59zFOrUwWbe9f2UfxI1JeNLHFTyk8DvjhVguCGg3agjo2b8+bSjK1+oDnm/G+cI8RgIoLlRyH
6rQsSOsoVLJPxSit1FkOaq55EXVWVwpojfRKJe6K35BAWae5Pp7vREQLN9dO1rP+5L3qcVd17n6i
sH4biNrNZVRLYO8szsWfBL2/Q4j1vhUVtcAUvgv2usYNbIl1peLfxdjHvPJD/8VuBxYWAHpOoWt5
IsaOvxVmuNP0xKkstao5TcgzacA7zLLBQAjWUKyaBFS/fJx5+g8/V9tiIL1JnFwwa5V9+NP4/lnv
gmUhUlsSjONwls+Gq5AuZwvnme3Kvm3kMYUx/IxO1ldk2Sg6Cu4W0ATsyI+dgOF4MglPfos3qwvl
xLUy4MgxHlwWqiiZbimcp/t2vfPewCTnc+VX2H95oFbpzSLv1Xb59s8pgg+IA/URFhw9nSuEH0Pl
0dOO2+kV0Hwb7g/6aSN2pC2Wz6S+3oIILgx5Rdbf/73yhwVf2y94U3RBaedHPJFAlxtOqE/bnlby
OGSA0yfjiXqB1R8YNb7hkU7f0NwLEzxQ4VKbCn/FHJx2HSxEG00WixOAPDlpdOl+wqFs1zQ3ln5t
8IZa4uHGyMJyfpXz1+aHEZlVEOCFGhiO1BPGVstYiXdxKXXIZ/bdoA5yl4pEtqih7wGU+FzpZ7IE
OerG+5unp94oaETxHBvOeTNj2KlYOMPqxBQdUyhCi+eK3bcZb43Q37OnjOsAZrKYtYKd2hOPfFUq
knp/g8nTTTJ/rz5hd8lS6aZqaB5TFU9HG9b7a5QpO+EUJOk/zY0Wd5yNthdYh/Bj9/4/ambfF4nc
b4brU4pydVbZl1uVfUMEHRn3mrCVVuLi/SI0BG9HzIGiYEsc+EE0YAYgCW/oTuycykex+X8iPLba
bvErL5fGtHCxhrVvlUaPvmPAIkue9XD/MOjUCxU1E9r2HpCmE2Tt80/JDt83utRvlFW4TxLzQmXt
9jZeopCCzPfcAqzTlexq4qdnGp5c8du4wgxgHBWfVjoU0NY2pmlfz4D+3ZFHmU9DvBYtikEQYP7l
7LebLQNHupQ83MgiZXPhcm89zBR/1ZAxVIYbtT5LgItMvbX4dAXbjdVdnGi1Nzn+cAFYrR1Rc2p6
4Dd8U2WpUgsfu51NzVbBDDqJt5orAI7QrijTPOEQDr5cqrPEJHsUacWIc691pGTHZZ0GI+cqg+/w
D620opUGiD7q/zryPMYD0IZIWBVkQJEtJdXqkR7RaMW8MIOlsz9FCJ6r6CuhQjiIEbyWwZ5ZbD+R
+kJIjqNzor75+czq18hwlbgKEql/fRGnFHzpe2kFJY+r1WuHztS2U5BaPpx2DZar1UtYa2ZgH7vc
KxaFgcb7LS6A1EflVlayG1Gn4vz2ZJRJkoEO/9EeaJ0i90nHxuvg12Xho/sPttKgZNVubzE9xsim
aKWAeDsF99YjtGNYmEGY7JDIEyqiOwj4W+XHoRdclnTQE6zmtp/0SaNdeZgOdEU87vMw5hFprTNE
+xzioC3HxqtFFCuviet83AQ9pJ9a2ZtvPBT8wx0JpzFW5tZPiWvZhBRi96ooaAfL30Qg9/Z/Hqre
AKrFhTcRAD8eKfZvtB5egS4pzcfgcENvbgTDCD0FnrtLAdMxwbuJhExxBjrqT9Mt3QnKlVse48yR
1uFcvtKISAx+Euel0NePxrI+ILH/MHxMrYo2etwTaQW9f0mi/AqrGYWo7OcsBflfu926ckELR5rG
voWm2TrZqT8mhycX0QgCqrwuBF//+lSscoEYUMBO0w4L9+r2HJprPgLPJ8It9LmGwqWGYtTdzh4r
Z5/N2Yse0ni2E/sGg/W/J1SaBGNzTLI6suCG9wZry1MtMgqMsHQLIFqtivqf18oimpcRviYYbTZh
lB6+JcfqY+px8Mh4eYVhbOFkM6DiVjFdXQXE349lZLaaFnBTagnBVz4SAZa2QeZAckGN0xnvdT0P
psZ7K9NcYH9Ka3d/btvdKvyjBAqRdBttz2+7Mejrro4gUCDQfkLqdhkYosdJTBECaVfDZ8vlSspe
HSCy9N65AkElWG9TMhZSXhn3ydVfFFGAp+mVPMtVuZSPN2LTLAzuUoUgwEf0pjr84f2Ry3Xs3Dy9
qDz50ed1HdjN9ZnxJbXHabmoSP1A1keA0wjIWmxgxJWK4j1hdcICVv/ELTYUwuKcashjBLM3uFyU
tKyVC8gKgr5eyT/HEwsYaO+4+gTWRCPfZDH7XC7MujNdWb3h4k9sKQqK52waVYjBCIVNNZ7VRLng
8BwRMuvBMc77pr9RY8/luGvvLWTo1mOolFbQWejTqbPfvrRo3XTkDbrJiedqbcIj0IHeRBkjQ4lE
+VkuA88z0R88aruSr3LWnuYfW60FE8SnQqY77eSmTFo+UhfYR6gmrfYYswqU6TwWzQeXF9vkyaU3
pUPiEpbx/WBDl1gP9xX2wr0fO0ZpnsELfr3dgCBXTfXJeAI8uqhFwIkW12kWu8AGSzgJB7MVMJSM
o76SIXGYpa7iIyqbUyuEois8LBJErEvSwipTbO1izgEjRr3gcNuJD5IOgl9RyYV/ytpfX45dwzVG
J1KeSk5slLbSmqpaP21L0qSgEOa9f9teD6j70pSkd//IYTcBihQuNUryTCtDYNNiA7EE5f4so+u6
hrw8rDAbwcrad/p4fXywHQFk9ZSTMd8W29pxqLXf8NvwdPp6haT3gs/GEF6QxFllityw3gRbbwkI
CiltltaCLVXFAojwP31/U1CfUzmibeUR4NAMEInnXq+fzvf/Bm/KdFyHvK4mboFX4DIG/0poEbO2
xcNMqhDOLm+RQSncKlDa2U6PYZWtoHxskHojEu8NeFz5dCd0yDbaXDMh95D1NeFzGeYB8r8i/V7f
lE4+KNnJQC3eFLB+oCBChMlF6o1PrJGjXCVieBn8au8wxJg4e10Rbbwr3D5RNt4VjlNym5SmqFJM
o+WErnMsJDIf5ELb20mEAZL3I542VKYHl0wKycEYGTiZpR+xESm2cUBTJhQZs5gy4WmQNnxkJGcy
s8oYr0M927nAheQ8TLvsahr/LoEXLzWJ3lTC7epCfAxfi2FJ+Ah9oSlharoxst+3j7O4i/bar2xr
dI849KLgz+MB8Z4MZGIylvaa2ChMnotQz7XoDDFPd77VrDheFsqYqvJbdIk5JrAi/32tbDQ8xO+4
iGUebeNV1giw1DFhY3SWJnAQbLSyHTBMGRS6WUBTLtZHp7yC3Ij64S8NH/C8sCUSl61QLRBwwEK/
O2vTF7orXLihH9vxVWVRVLpjRthlIwJwEYA4E8PkP/g2PesjHci7hb3EwHN21XkImOCeViS3LEd+
EZps/4LeJqEIrPXt+opkLUEWXCTlg0ZtQtmnMufJsgvwDEt+336XwgwyP2IDZAGMBOO2QpdMOISJ
iq1D5OuWnojrNmXq+71X5C8twUQiNOWI6cZOZAm62+HyeAbjAAm5OLU5m3dhQLErO+e0Y7DGQSnd
WPgyW8lw7UbiBXIL14rC7dqLXIRIRpQ8iFRiZaWeer605UFjfwGAs/GlozCX38fZpfTukVaoS0jT
lGjt0//YafEQGlzSblzGQDBKXgKGwRUtn1/DLYDSKQkyF5IEbsrDTRAiDzinJKTSaGwmR1mKjsFW
xZuT1pzkMUcQEX3ADJPq94sBY9pKTp4nmUjbKKGq0l6KcnyAycY8rlsQU0FwgNh0/D5fS83eJ/Z8
Q7w0ljAAKu4SUOzemCJqBnN/+s7Nbwir9I/HGfY0Dr3K5ShA/F5isBYUMPXAfLYz/nv2BAz4KB82
c1rcSYTfgY2RozlfkDP5RGln2e22RSbsKzx5CYfvRKAB9vTbFlKmp+72bQ9+nZ+PUwLSWMdSO88T
F8ySeQHi+YB62wFF+uxsUNXHSDF931s96ADQ9MMGnUpugaVnBM4/ua41XM3zN1bK0iJcvqW0vBH9
WDMx0oFVcVpmRqyugtZ6JBdu8dL1DKrq66U0CouNRUjItbtVEn9jV0OcEbObHetJzPUEFlUAaLPo
bfflRj7A9VicTdZavOvRFRrPAhF6evO6h0PKJwDsiYn+iE+MXaURHnM7QCfw3GSFLgVBHHm7kzyb
D9b8ABLuCiRf3Xa5jHrXCFkV8DOK7BtZzwaZKBT2GQON9WXxRAtnoJa1T5dthkj4hTvIdYT4R7HW
iPQ8mAZWoRlbuRPIQIbHLFT47vMbDO/avOREd13Jb35711oJIA9EWG3grq3FR8X2zhB5a37tMPKH
dsdr5W57vnw4FInBtJrru12LiJkH6SBXJY0dAJSIYFDGJZhwSJlS/jc3Cr2mgzQrYZ8nSL/HTogn
vwU5wJyTswErHaL5/gnxm6l1eGTSuUQALwbw2KkC5XDtCnC0GJTXvRhQY/PoyChlo/KkwV6iUzI8
QSim3AYqy/KNDJn6RbBVU8D/JhLbt/YoughBIVVHGkkB5A9d3sp2qxUOdNqY18JPd/3BEUgJ9Sy+
YI+f+EWItq44B2xduN4L3mcbGEStWn+jvTm7RdS1iYEbL+xJH9trVBmeh/sN/aYhElBNRAgI65pj
zFXV5oYJaKrxLar88Ksl3zM93xsr+MN//h+WSfwKhJfxHgvT9mUNWAGB4szZRwQhFfOd93sy9lYj
d6LMa6zM0ishSvLXIwcZxqvtuIpIUkqlXYJqNNMfqbiIf5H5sBv6GoG7RYET27tupjFdTeFC2RFx
7cp6Z9thPqSE+1h1U2ebhqSl7MGvoth6byf6pCVNQHPJC3UbcPcNfmm7soupP7+lcI+X3Og88JGH
4qlm8gQs/5srgq7F8NR357rn3lCcB3QaKwk3MrLVwpdy1echc7hHpo7gD4Dkf0mt6nugJ5xikCKa
+RpOtgn9ouI6pS1C3LDHgsBg8oAiyBmqLu/TH9Od1Srrt0zzrNDrROMHz1FU6WvuAb8V4rrOkU9H
0hMhw7WCR7foExuvyTmHOtfif1TfVEZM/0W4KIGvO8bf3yVwAb0wyyXmvgsg1ikaNRBfKGxxrv2N
0c8gB/iKlcj/VVmaqpFkPZsjtEMPEtELtsxrbmYVjwBVaXXe9sAJ9mX8KU+/2d4I/SQK4Uf1CXHO
54p+dYzMWj/82CmJMiBYoCbsMpzpmnthkl0U8sHvsiTjn+PpEh7SGJFI7K/RGJHVE2xIEpcknYuj
WXCMa6uTADRd4gR5CqJW6iUtNOUQEhC75KDW7+cZhsn41570LBJkjSqlYrPdkPAB9pfvboT/uS6E
galBh6O0fmGoEYEL/M5a1CF9cJgdwLo6mfQqV1vZeVt9htNbJ58EEfhJ6xV5HM3ygfpsX4mFLnH0
Z8iJkGa82POs+ajW/6ujx+lrAhj+/XA+F7qgjADBeXJW/CQ6ZInawxVjpW4QrmeRy+i2l2XJBtjw
7CKkqBOplAsSlD8PcplNvCIeiu5Bfvo2D6jNPn0dcM7rOsJ0m8gz/Jy+TpafYdZ6xqnwmCD2TEup
t4n5KkLA9Q4BYpfB9Z7D55HhV0Yv5DUHbHRz68UwrMj23sUjT+gGr+ZIOjsW3q0fF6wWy8C2Xza5
d3PHPK8LRwDJcsUbLeI2J9k4xUXNslAVJ/Z9Rg9LMfIq/S+kSDK6Itq2nufMZL/GiqYH1jpvqBmz
Dx1DHHyu+kfXMjp+7cGswAnVe4GyicScIeewvUZ8pzxLl2PrACRhBLigXWba4hn6nUOIVg3+w9I7
BnkoIp8CXZJUGbRBwCSRodawJEhobyY0z7PIhNjzjxpzilOcZt7wyRNNYdJTKXgMpXnwp8Mu1bqS
ylHG7XVFrhBZLwNb6CSZnepSETBOgYZ4Kw9PF80jgErI9xffs42JMEFt1YLV85111anY5cTjUz61
qBiva4qfAWosjMMoBcw4Sp11WAKvGZlyH/lJg92Zt2LnzO8uo3I0N5UWnT0AfZvi/CviYOXKZX36
z0jlEZMr/mZrPWqIviDG1rAqKFIMtiVkGgr49bvaUdi/TKxMgtHcX9vnaWfyzdQBSaWfZvVjEvKe
vaZ+YARk94eVP1rPztEJu8tPWYbZpJqH+OoSj8BNhwUiY5IKKVGGpVprdjN8Q/kwBufNnXeHCTu6
6H0RrFPnR9p3NPE9dI7iLDOqnIRO+iLpqmVj+JdNlN4uFPqvAMnBc3Rsu6ypP0A5ag4hULCDGYdT
N0wnebuE+c/viHWIuCfVmxTFzoePGtjXXho0/5lZwrpc0EhCpgPx3b8fMcNxbKJh1kgQVQmy5G0t
zXcl5lIbp9ZhQGaQ2ppRPL38VCD6b0mt4HHFvbFQPCf0+Jy49EuKFxTldKF5Ay6C/jwNH7/XrK56
qTn2NM2mqGcqONu/GJShO0XhyvWrIbxgTFLzPgdT8wYvgPcv6a3pqvwC3UfUSeH1DPl9Qeidcvih
ngyAJyakMsYE7N/nfR0tdvM5v56FqPOscFZF80M4wRRuchDQeer4DnO5q8d0Xwf1o4XCEqHrDODB
+nGLYwHcb2yR25LtxeEXjuLOreoJimsm2PdEWVb9p710dcjJMAuC2oSbEmyZQURkizK/7Byb2KX3
7yhm9mYWRIO/hbbox5v70dWBC/k2TQ3ajK7hn3DoyXYueOPQ2IxliyO3znhmrHPAAOWo6EKFOBEH
gY8Y4XqbL1BF9NPmHNaLlVpcRqLVkKfJ6X0Q/MTZrvIJMbvQhIufcfc1/KxfFozRWLlUBrL5i9Ch
stUyZ5wVkA+/89Fynt7XXp9RCaDo5D2Kq4yE4w2fxALrzmVxN5Pl2L63D/q8NAUpBCriQ6qEans6
xjB3QES4Dc8GNw282VmmWlIJD46yf2DXCsOnu6MUviSE2q3wuhhHKPuLAhJSM2PItIZSzvhGJuqP
1aT3deTu6AlB+1ofFBwcqa2ABJFvx3DDYLa9zuqtPs29LgggVeKrNvW8hqCTapV7YUvWgK0dhabD
eJS3e4HqcP+pL3OtcLZvfqCI+0xnfMx1dmnFXJjTg7PAsPXNTStA9Krrx6jAfwLUZZZWfdfiRJES
jsCaJMkRMMaesmifzYmvq2aWzxTd8NKjM5Mzw+EkhdyX+n2CvFhHGU/ipuLfKJsd3MgJA8TOoyS7
a6yiBbWShsz7nCjK7lJhbKtIVSEf378yKCY9QtnTZmDX7chCikd5QY0DdcV6eLuZk6+FsqyWJnVK
B0WhaFtS2jBIgXY+TCeii9z4ZpN/b2JzQ9PJ5j4gZmAUb/aRDJNvv5DBgnIlZKNnsoi/smqGvMBW
y1dDxAsS8KljF5K2zhDjm3J52Eu7Ye4zp0R6bPHY7u+k6cCkC0aOMOOtH3jp0OlTdRM9cXziN+Md
ArtaTy+HC+wrBXwwhjXwDuroGNU9GwpTnXBQGdwIzoUt5QUMs8jX0M/ejKBxvaim7lXojep+oXb/
+8IArVgx3/Nl0bkj9z34My1de8noEnD8wwEc5vD+sNP7QWQm9w4xg/1xRiExvSAFkEbHXura8sDL
LxlyRzu+MWKFqfBgjFqmtRAaEg5UwAWWLWE9Zci0o/gOoA6+UDu8FgX3yNslAIqTJt/0DPs76pSN
IcvOX5OZ/E48LJSBhkOADVx95PF8kK4CHJM86u/QcPzUv07z51BHMoCaC3FUsATvY1ihPpnad9ti
+uARGSj1fRrJdJLFR9Nz/xvmynBs1SiUapFpKOc8Fe/S5cXLCeidbxQA3VuHNo2DxdoqFFPu3QsS
woY0djyG+0u+cGnkihOedPlDyCe4h6YzhNbfH6Gl18HJPxD3y8U+bpO3Vee2wFwiBzYquWeAIatn
BlqvsNma6ZkTgtiSLBeNiJdAyUFbKF0LDaCIe+jkfODKORtnbAxyOcXH/4s8G6j5OtNJA/Io3hAZ
ZpjvYXMAuxPhDeTd1o5DOBUgWIn1gzpm5PeHEZTgCoLZbDNXuw1oS1YPHmpilN65KpHxbvufPfEn
sWBWFbPZvxxx7y8fKwy21cIefd2Zqa2Dqw4X7EHr1FQORDGDc0JSUS2Atb+8XczknoIrsZg7HOQ2
GBC8zJQ5msVosO0xNVNzV1vp1wHH/KlnAHm/86R0X8G5FUijHVnMShjZVHqLa/7JAUSJ8i6JerGr
eKL/3x/1l95exRCQeQDlr4YLA6XXp9nkbqm/LbsXrBcNXYJ/Yj1O5W86dtSAG9CTzCkdf5NxB12N
Ujo+gFTBn0kSAzYEZiFdUMFkGwd3U+2gv5Xp3wd4FkwO6IRrg1YnZpfImB1f7kYY0/3N6L04L6Zz
h0fVdAZhKH3FxMhy16XyZvUMBbwnNjTfm3XENi9IC/R90hHVZ9LkiKZlxUubyd6W6MGQ5rp+ZQKX
aPN26K4jDBXfkgCexegVifNuTtgGsHw3npr+3IFuOm/4S9O+kg4/xw7qYwgB6l+Dn9AEG7qS1X6B
3kdzhcuKKw4BP6Q395wUuP2pKZeV7r2Rmyh7ja8o+nH8e4kbd3RU7NOCJl+ao05tiObdwLkkJngn
jPidtkduPkQdKWNyHNNDSOdgX0gvGsMafN1aLGl75/uFjfPM/kq1yOQeif5aspUe1bMs5a73S4C3
Z6vesFveTJ8y4mXrhiwDzqoDEoFcHAY4R7gifCre3Balboua7ZUazYJu2w4TzL+tBy1Ur/I3HaxT
cuvyLgdX8r7MWTaSW7ZltittCJQcExAxKaiaJAdXr4o9VYmXDFkxd3BVZVohu2uUHn1G4YwmLZXR
eblHl54EaabTAzH7YRusBfERKUN7qaQUrkKUi8dfPXOhWgG3JneLAvMaUE+MOjLvSsh5h8kk+X0s
1M27zgfvoExvkG5Quc+k/yJsKSQ4M38F+FqqEkMUMyw8u10O4mmwejqmKmN/vy2O7BMuxc1jZ/xl
YtLnSZdtCpxYrQzYlI0wd+5RQi6UslQNRBcSaR1naU+C7wjuXbfhrkordHX31+jUnNUz4PtSzqwB
8bZZnC5CUa+xw4mwFt3TM2iustulCzQWarMDoxPwzI3Z57BXdGihaWZA+y5u/N/KVvOntN6DWen/
YPlj+EwG1mRhBxhq9HE4sMSTZd2t0GE9berRBd8wRYwThuxQUAlYoWR6YLslbLs5eIslHjfaulxE
rE1+e3/26JICWX4P+Bgt5ayEN7sSouhlrvl0h7Ibv0BMLSeHJexSljvFQjAHSQAvZUko6+TDiXmJ
g5hNuoEYZw1r3rIlAYMh7G/cxe676+h+7fEEwX53ovqd2J94R3bAcyp+VpL2dbo4XLyUFMfF57ft
w9YK7P3pXIKt8b2He58167AMc2ln7uxMfmAP8Au1LBuMf6Fm5YCz8yHm0T3cH2ufbbj/+ovQoUDR
/7SUgwY87Zzr4+BJq1a9hudT3MFPssLYaT4Y/YHOawCtQBQnxbuQI750aC6dzCaelZJ+hQ3O8RFk
SGwB4AEz2+u1TkBtukXH7KK0vZAl+Ptb0e6RtbQ/ssPAwQD/Y/l2GnMjXFVcWOeO+5ZZybyfOy6Z
Nc0VeX9RZpnzLyRD959nQ4WlrqKhjDD9f/SLk1REUW0BUk7EMcxLqf8u+0oJsIoQ4l1ZF4tE6b71
uTNDm7IjOBm5IzF62ibv5mLWy80NuGwf/4+q6LQxb5gySv8qhyYfxHAIO715hSb8JHZKPzOqPcEK
CLEJABpOzCsmVru54sqgJ3tIvGuFS8yNSXWCrtpwB+lhOIQ+t4vhkuho5pofzw+jXZ+gooKscRyQ
6s7fqPgIYt7bhjf96wEgeVBJ7giaT4Ncvq97DTCXz9hQNScN+6iyj9ZYTLQ6YKZ3YAjMdTDJShpQ
6kKDoxNUQlD6Ic4HWu7/G4i14YsaVjzPWoFUfRuDT3/zaT0dXPHekn0XDPnGGYaeCm/5IviCcD1F
B8uJPxDZx9J684Xb84aVlbrUiznhQLY9FpMAscBFbx+MnK2aLmPaGjN/r/dl100y4BlLL8m5pxed
kUkpmx8WBZy2x93LOXI/EysQbjfa/AnrlnmozOgTEY7uE3wey5cACzLVIPzcHwi7GJj8IBKFbQhO
Z1ah5n+BzXo4w6m9+AeJZGKxkS+iATPjQCeKwlqOIkrvZYXTraTKxD9IJ2cx4QHqeDWiXbqVH7j/
0Bz3FVkaTKPMbjHM8UeiIHVIt5gkP/OmXr6wqSZPpLNGLykYJC2/1AcV9+P9htf9UuYalDv1ZqAd
6RMyzpVBsEp5a0DtkVq40PdRf2rWtaOcW9tRdPYPH1EYkZR7dq2pU9TXxH8pu1p+k56U0oUDUJ6s
1e6hY83vZXmd0GUBqdLaAwaEDVHmlt8c+CeJnhR2OXRA7NfN02v6sgc5Bm4Cas2aamEaXhwslMz0
NyVH/xJl+JrcSzldGTJ362DyR44zTDc0prpx/WADFeuUwisa4zKwqGFIDlu7gYQTdWI1JMgqf8jo
q3uPEaylD/wCft8SrkBtKZ3LskwboMPuU3uFDCzVDtX13IY9sU7U3Y24K15nli7GCrwtOk+njk+y
vD/EVQH+hJyjNP6+ZmvnA2Npt9bqoIY/FdEL5riUlKo2QmKpfJvGzdJRqAqhn7g4N9dd891alGcv
cMIk3soyR+dvX5oxzhOIdYt+Y5sne+mizSc+Xkr348IFbhnM3jSzHkXIXN/dBbGgMTr5Sr6Zmi7Q
QkmOD+FwA4hjkC5aC+RORAWTFaBiOcM2PE8F4OvZpWDDhJnA5MG8/agG0eMvJQcfkaNW8txfOWqT
ue+Pfw5e+HGz3shDt8+6VhIpJgpudre9AtSIAjeckIxArxODLblSWp1+eViwDd1MRPRimfjhEcOU
I+x+wiMx9+UpIbkv5WxIRBszNdFTg9V7ZbC3a+G9oWG+It7oDhsByvGmBM2r5cOP/S8er/17kVZb
Ahay8Hri1+Lmb3rLV/vxIvr+WekFPcErEPgBEl6aZSNVGgVpeBVtJHGU6bxTs60sYZHBM14cR7d1
3pBXkw1+ea3UHd+ot+DbEU7OseQm/8CVU9e7Gi035/lt1KZL0JsikLz+A93p7j+9kn5DdVAbv7P1
JC8P9JDG9Nd+iaJ9+gnl3DeMtBibHETHM17eqbadE3KOPg2P37q3i2MLjUmZ4t5Mhkt3Y4/BhiPV
t3/w4nP9YodoqWFrRyPoWo7f42xtKBj4KJ38W9hd60z8uY6N68GYbizjRFuQrVBex3KSj+ISl+Wa
FbjchWBfiUdzapEu1uHj6OhN6O8sBYSbLyQMJJU9XS+rBcSICMLKyNspJyoalabQQ2FYP2SaOXQE
QLsLzQw/BAfhPZ1gOR08ZK73otAr8OHeu6XKFtADZkE70uz47IUDTnoaeHvncwbdc3UCdXNZSWUe
Gohs0xi1OG3NUPpSthhpEmYFB+27PsQOMzKfa7y/qgECEvsdT9bfIJsalAW0+kr9e0TieosBQD89
faaVVpC5mg/eToqInMF3fPLFkmQBkgie70CMzrxaAmUnKOSc3ZcWmcogrES3FTRpfMgMZa9gXRbt
GAxMsJJmmGSFsgaDvMIiToq/kLkiL4UpOAdjzEvUs1w7jj5XbHmM3npixrqKiaUowMR9QcxEpVXN
oFE5C1CMqNdJNsZxDRiOVXbaBiiRWIwjDxS2jL7Y5v9yHCTOwD/RL9f4rfiGkKa+2CHIxNjxuVZ/
KKajRVmHGUue/MEMHdYfvM1cxcZXqTnv7i/Pos+19qN0uE43Q/VNseNTQwZt4ARuNKO8AxkHHn68
iqATcYU+G5PwYqa1N0tL6pulkLKdEOMINsgMv5lDUgpeuIZtwcomi+BtzNfkPwo9myzT5MKtnDVR
p1iTrcCXdp9Fu6C+hlB0UY7wkEIY29RKcX8eciEtSx16z1WsZDCKHvgjPKRPB8FRt0GMWoK4jyaQ
DKt3aIxEhtdBGjtJffG5FunYhegne6lb+/YbTwU5O6D2mmdNXg8cByqPv0GoO9XUF8EUJ0FtEd0E
D6ZjhInnqu6lHf1eqPsqXxJ0Ux2dEhp1fy8xBB6AZR+dfX9PrlzyWwqXsGhLSXZ5aT7XRN3ClGNN
9MXt4mUcyuXzohYRAFi8jPRhAVwf0GMrRN+M90jL2oKp0ZQJvx3fDIwWnk2YfSzBPF5TgKv5pA7y
YlsUyTNuoXaRpEapAcgd+40fxCBSTlKzcsACbi2sTlm8/COxj5QgAtbNBWqUKb6UE23lLZdYRobJ
Kh2ihmyztvYBW0olDS8Y78poYgREG4K6LvPPkZPKe7799H9DnI+reYghmhUh1XpI6iyAJIaYhZBG
516boMXlw9xnILRY8GqBnccYQ6QuHkX14iUwUzRvi/pruWH1hUD3CU+CTZGEU7Z4s461eAslMU3m
EDxL7xtB07lKmGE8hf9Vopa7lCwcIOfuK2bHkHaCjSTzsk8nbmchRo6bifFxmOd4XfJZBxcs/gqo
T17l1PN4CQ66M55Dsw1qBiJL0i1xKCu2r4/C/wClSsyFuPcmtIJGN6szdGx4savIPhyigETFH22K
xNJJFdwFt6AIPDgexoLKBRqKKE5NzqwpBNJhWg1ABmlaQeRMbM7VXor/5sLqiOjMuNg7RRnYG56B
xv29+gkOXpEnyTakqUlY5oOPEnKo4B4ECOgSoe/FfMjJiXePJnwFKa0i0NYo0juM6tl83lJkjUjl
HvaQz9bx824MFKcw9QNmwNxQZRE04t/GBLQOQP9Xr97oN92QfgIFpfNauJnJeMkqc2Hm1kBI4C02
/2WhC4WtoqfdkrHlJUf2fGW2ssuqwRK1bFzhWmbqo99zc93QP0OcPA2OKvGxEgfbqp4sEUW2B/vW
V529lCPh/xMM8M6jr3t8u2lbu/Ug6SJetWn+CVA46nZUev+sfhY/ah9/a7Y0nOLkDw7hTCyupWJo
qi4OFAsBE1+bCvEO68lE6tTra4M9BsQlSJTFbrVNqzHzPQV9snKbSplB2DpVchF5nXTjLCbUCv+C
q0xtNQqjBlkgXpeyCuuKmrHThM1emBkVNgpd2oqqRDSuy4DMAYgHGzwjoyCyMu8nzJsDceTVS1OP
4M29Wt8LqX4CHyANktjYOwypaf3Q+jEXbTkrC5BljPWrYm3gmAx4L1cq7E81e4Iwe/nI9nc/rgBY
XnysAS9kHZRL4YO18lHXsttjdMnyuyk93ZBoGSzw0qQfiszvQUnSnVUyeoFz1YaKdEtjeeXGRD3R
ACtaDpTAtFkz1CcVD8pXlhZ+hLo2srHl9V90UTjprlqg9c2zJ3EJdMg9BQ5CUAl0eNCv6lin2CCl
xRZIr2rqGQeQWCkiFAKE6MyKh/lU8yyafSeX28kMJUmM4cpcsLs+7ssSqEEifVI0fIWUpLTqiJOa
9GDVxVZ9obrjELeW/qSMvS8W7DxY6PXGxYvSg0VSY7l/l0JdOIfNHfiMjIKAusuuz03IIIGB0otv
PsnpTghyWeKwmTaOyIXpVAw0wdQqFdLJ09muyKFLJ8n9L4jYEmLCMERQhQFmYf2AOh1amXgMyk61
7dswPguz8/Q5oYSN7IsvXnAyeJZibAgiBOAyieAWLhbtJ4Q5rSDyDvgqU8hJ3PPYZ4dS+wB1WZuQ
97vO1QJAQx6uFMK0qCcE56NLX56gykhFMoz/xJFo0MYTVhuXZADQbC7WTJwdZxAFJVlyIDs6n10m
FTpE3ALx/8yshgZ70vvK6VbR6oAik5SP2oKWc9fvLc8mhsaeI+3n16zEEc38FLuLmWrNDG7k3YSV
qd3zyBcNgOsJgA9oDvURVr3x0aQyuqfB95XV3OtK7H1YciIQrekWGtw1+iaeIVhiGrSsXSoiG8RQ
yOTv3A8Tp8ENi01YZ4odJGM5ATY9HkCGwobTl7zEuLVh+VDaBLqoPkoZg85nSRHw9R49ocOMN/Ww
MVZ7+DfYciQS+OygUN4IoL5bEvZJCElL1F11t8goUFdOU7kjQNob8ZqNXdlx06wa/mayvf2vGbIM
xy2snNdKHYDhe8NoF1n4o24RA/QbqX6hJLfw/23D9LkalCsERO8zvJlfTNy2XNdF7YGkPdwO4PLW
sASvoz7/waetkyXD8KfR3GDS9QgrYDIpXs9pefRKU9nucIc7lmkA1av/J2SuczZiFdNEV1a9QvUW
Mz9lP/Ck+aC8+2C4umNiOqbXuCuKdKYyAviLDIn27lvY4BlNBJAIwCWgB8TmObvgZYLy6Ap0mZo3
X2bKWV1aNjpdOJGOb+v8YBwm5sMTWTEzZaiy9Qq0/o0s8decfjutO98w4BULBIKWPyPtViN9fl3F
apGuiJAITX7mvrNvmrFUmf0NgNWsyT18X5gSxgrP4Rwi+Nj3q60D1fQCMonl77WDM9NDgbZ8Tro2
YjT2wyYO6w3CKFw8S9L5euFxFg0uZsW1+o2sfWdVjOQ3RMeaJGNxBmxjpi86IUdojH4w7Ypzjyz3
bUNdiRU8MhJ/vew+88Atvhs2RJXsX9FoJpsimiEnK+1wh06UiGizkmpMu+5X2FmGLRwNIHu2l1f7
l08c9SVPPU001NoAoikXa8ii2LMTfC0YU8FyQiH0hydrGexminYDV3KmfwT1ew+HJXrPcS1lDu8N
cLy5hx2I95+FXoL1LRmXSH0VMPLvon2cY3+PdWCxFUiXN/0gY3p7o1OAjwDNTwnDbMSYVcKjpDKW
T3EdAJnQl1WjpmR5hoB/xXH2Z4Iee8KJvOGGyz6v9OGeKELEyMTe7UwjrMULHNZwVihQBscoARq9
URa6UodqUENMl+R60aLYx6VGRur7d0aEmGP3fLbVYRyagh+lF0hluBhZFhSdVKw7e1dUYFTf7iXh
MsO9M1zcxVKIIpMgMbjzVVSSYlFys9eFVjXtLKFbEJaRfz2DIM1wXlN3u9MZSVaJu1NCAecPxI8Q
pvqh9ZZUjj7fYelnFSgPBxVgtyWtidKVRF4wx4KsOC4fdmiYFNfHwbbiUCHZbfVB/af72pJBHNnA
6rt4Z+VKQv9a1HVievYC2oDG/bDVVld6wpcyukuvh7WinAj7BnBmLc2y0M8e8vqTt5Sm0doRkS8a
sICVYVLaF26+VL5RCPZmpMr2hqIF9Bbkk30+sxtU3wfhHrIczcJ+D3G/XMmKGlkyXYmFoXCEI5s2
xeu3e61s2oLQ/nIzbhpxsPH8p0DFVai5TUwwGLLLtQeXrL6GyNF6w2G3e8AQ7/vY59xiJxTbtdAY
P5R4Vy5Elv1ncwqwogAEXObj4K1oVL3ATpG7S5iujHfcnX55cCU/TpUXbOKopmf1l//CXHh+OrxJ
XSp1sQ7ium1IUwMu62lj1KWSoC/+yWeE2aXJ7c5wmqIzke760RYPfQ/1LD8M4k4K1ZWiPs6R92ik
AtmO6AL7Lnm8jXHOF+29AzlQiahF6BPlrunjK9hSkAEY0vCG/KWLpYOPxuWAg9skLPBs3e5Oowsw
LkUTNwyU9JRriSzEN/yRR+/TrW7UbndoLFQnyZFkfnIftj4AKuHBWCFYUQJtbZX10zcSCVKpPztP
r1v78vBSpq3FD7bzN8ySordVcIL59QIM82r48VDZ3JuBdUzWJ9NmNI7UTKf8OFzfWz4DZp1KOmOb
+sq5EJLvoGxoo5adqU0bMmXbKIti0WI82MBAQNdWXrVKyD0aZvKTCYrKq3IJ3IOYlohMBg7ATnCz
B0ikZ+VbOHa2a0PruwZ5mN1agUEf8xFdwQ/rYZ8C0eRtwL6ub/nqBG8iX22m+GXHvUsOEXKrtu2G
xQDt3LDXSDyHMoaWV3AYxU31w2xgmA0P+fn0FERYwTxGHfMWu/Jz5r5B1+q4RLfgKwECg1vdRRGS
Y6s8h/OoEsutowE2YyaLVNYbbPGa7aLzKxpZOQH9P26vDvFoV4VjwIO9GM3np3Frc1rDA2kbI49b
pOA9sFyLgjZExMT48AwdM4jKSEiRdnyf7uF2WZh/PZ0FVXRVGTAb9KKXloe56bMxfBos6t2B0B+G
oqQmqxivONC3SZPGOekaLlk/CtPrTOP8pEl53z660HUsiG81pZM90BrYyCQPftVVI+Gnt1+Go6rz
X7K+hFULpCUf+TtyexxVkfSbu0WGg890xQk7+AGOTou+Qj6KKyHh6QXI9MEAd8cKxDC1tHhB7pLT
9KQhqgnc9IKK4AqpCHsSsgIdUVRA5ayBzlpaSQV1mskz50atKlnEpeTJcc51WbMUyxfboLTIVs4d
WfOWruZlDCvFKkKXmo8XB7KNG1lL7mM9q7ALwgIpIXNkCqJ8/PPLZNJ2V4DZJuH5n3+0r+YUJOdD
b4LZHVD1IB5km4xl/W9wTb+bjS32HO0f8NiM1PrbaIr7e4e2AO0GWlWcBo5aJFlGiqufgEJcPHUl
k3WCU7fh1/jGW1jpp0dOmzdbqCGMtbhPVU8Eg50Ulaxhaw5t8KVAKMuqe/akwFJS4OIaZP0bud2i
8BDP9/gfGZ8d3FDe0JD72tuEBfHJUnmIUjA3lXJ42AQ1xqjNZOwTRazqHnDxd7qFl2UUgXRpaAto
eGPzerVPPpTVuH9AswRWzXn4d1aaSKZMLpeVh5+UMI0t5orF7PLAhtk2wzkoixYxbx8qmi4EThc1
7nsOoixF9nxYdhQx7owodwXwQbrTSsczoyErf1lU2tv208oPLqSgaUulyJQLxOGzuOusuYImGQcH
Axnw7GxeV37aXRHkjm2XGqSofLY73UvTdcEnipXOCftteT491oGJv8khCFf1nSL4QDB+M4HeWteH
Tu+2tbrwq0HwOyhq7XDQSk43aDNHRbVdXdA85lDe8X+2/xL5kAGm7ZUPTIQ4XyV3xTed7ty/cBaY
KV5BUuABZGhZ8exd+AxrPr226zPnxfzajzN+HWSwGmYLfEMSVOM11IqegsfBaVBOdFFQXgHZUcl7
k/EuR3SI8ze3yORAnJWi056wZo7PubHy8I/frIUx0Wji2D5jg5ezi9WIePQ2cechVcga9tAJgw3P
qMn1nKHa5AXMFxsIwHdpgtg1N9YV2WdtscWTdOC0AZyYmC2zjBd3V0Vq+7jo5HwEgf9WnPPWTT8x
Xlh7O9kPeiZt0sMW+pG1leLPDSa/Pva6V2AP8fr4TdhhLNz5+nMs6d2/n0613yYoUl9piJOkZ73T
hMAjS/IZwqSLd9UxQTvrRmtrvBrUcHaJT0b645jD7695Ejz+yS+cwyroBuwCq7NW9Cq1fS/ischM
U7RgmzBu93d99v3rga4C74ejXNK2YnuLK3ZBQ+hKlUaxKhuocCC+P3cddntxBPz113NdJW4uoAhK
4+fdJVU/kfkrohott+XcNZ4jH4wD7MNVVrq11JTRsvfNjidWy51zz2/5p8a0PukxRILllLoXVk+A
5icHYSYarQ19iUQ1Xi2ymcLFS7O2XDwWK7UpJfEbQuAd7XGHuItDbaje1sGvzanGpNQUlITx+wfk
wkMcqgd/Y2ZDuiCdKoOuNLcJ9hgnxPnHHk5LnLG49XW4mUxtYQJjIFU4YmlZrv5TYLTa6eJ9eI/8
ZXSatJxzSvNo+41KB3T5w2htOLj7lWgNwxGegs/M0FzjvjoF2HKt6qtTPuUsomT86SKrwhQcboto
mI128iixXPWYTb0VZRupawU6Ui+Ui6du+IvdUpTpLRGbEE+t2bxrYkU4cH4YQhcf4TCK3oPJ/y64
w0sRdAm2io+YVbq2Vrkhw/gbJtx/Fnp9T0UJ3mSTizRIYJr/NMMTf9wtjxaY/0NkOfskVknVj56v
ktLRm8mcmuFHCyKL9mhPaNgO303Z9ttell6tbyZXwEG0y5lAEkCluLjP66I2a20DSgxJ5PgjBgXe
5VpJEWslUd3xTc142WpPrmNlXxkuburgMx5Ne+5/J/TYNWMLjjLIDBQ+TbJBer3Smvwwr0MCpetI
YTiqvL8Woj5pnkK4PhweUf8RFvP0XtHKoE5l7ORIYOvS63ulYjnavJS/PQwk4c9YtbQcJMO1iTrT
3yVcBQFl3VjrTWfVwEHKe6HZSEUUxoegOu/7JBdP786yWAtDATrIhFG3CCTQVLe3XBmm2/ilzEoK
W5Rtu7Ml0c7U6H5pU+vZqxfnAN4H5M0A90GUM8s19HR5dumnC/wJd7eTJHkUXsIgcgzT7bT/Bsf6
GCh4+3AIUdq0DBbsrPvbUHYV/SR/6/qTp/RaAOypi9niJSEkgH5KjO7wtxUIuYoA1mW12msR5N4r
Dc3msyARuKbFoLbAp24dAqXl0eWvkwkCX/S863imMaPlsUKt3+8w5x4a8wg5X+5CWKsck7pOREbT
844WawTh1X9osuHF1ryi2mZrwTwwMbKHTXQypoKab6xnZOFDpLaZvZI7OnvHGAWZ4Iq83aZR1ALn
3a/tfOPgnpKgo7qwIbqFDz3KVNoonebMt1Jtv2c3btRanBNkvJrcyMQ1t6UswPp2RRzt0TqBTrQe
EyrsvGcRAo6yBI9MI4G1i3eoRftjP4RV/gtyT97BXBYyIxe+39sNqG+dzsBAY9GES2Mz7q6Crkk2
f6YWaFDSx1+uMppKHk1wgZbhzYOtviJA0Zq4u7kEuwTEnGsSF6aHglODIFTBHlotR4Hq7yM7cGjk
SG8tAKmge65F1bWonxOTlGKpvYFzdsokW443JGBToj7WNfsYLG4+tmlx0joy7HlgcnHH2X7DELO6
BbtzSCLgVrklw0atQLvmhhmHtEzU8HUhVogx+NUwVAMbFE4q8gDattqiFix0p3qvd0p19dpx8uto
FSOOrqpUphDD/gPAOkME+nSfZe7Y81mWhi8bka3jxTKsJ2P2dcxX2zk1b2pXPQxwcTLQQFTLcgsE
JyfTzl0j/p+zub9BEyn1bL5RS8fiYl5U5AyjK24H8cv5QtahEk1XSCMmBppyg2ZmYNLmvwxCNLv4
Sueix2gWnLvGOvsz+AZI5rG7VgxwncGa0KazSQB2WW6OBujaBeDAyPXH3fXfhZ0gYdtNaoj9mGud
xYMm/hW22EGrGpbhpXifOUVpNLcs/5YDaw7UM8B59InZtsAOIFqZ2gCzmXhOH864vDfE7VvVhHaS
kSTve63OUpW7LwYGXHBBs//cf7U3akR9yvlQVQ3KVa3Nx/2FckYapuqS97sLqf7zdXtqHKVp51sg
c7kP2wSaDtW2Q90qhCv/aIXGKNfcbw+gcsTGkHa1r5AtK3CFW77/HTTabGt+pNCVxqgmNtS4Hk8Z
oyzLh4RqMFcHp/p1boBRkos6o4CuOoRgMriQrP6k4/NDONU2FDzgK24CJ6Urn8wg6ucxnUl1LgOd
ICOjg/zjNAP7eGQQ2/0qb7UVc0mhmFi2Ckzmzxm/dJM6wvg2399QvYP9zemzWucWpTDBo1Cnmn+J
dkQvcDGZHsz7O6+NtLVPl375Tn/hew6FSRlQkH6P8NTg8RSSL4SNfMc4ka6OrOnwAlID9U8ZP3BR
DfAW5VDouZwwZVIRUPACzXz54Xf9qpxLElUppSsUEFrgVc+VnvPRxpIhGM7Gh+XDrT9m7Od+r1f7
tqVcRYGDyagGCAN6O9Ys6H+X9Ax3TMQZ9zroNzomzd2NRnDs2SgdIfqO9hMOiMUCjy2pei0Xtk3g
OpJPZnWktdWkLEkNC9Ffg1+G8QUiGxjIlq3l1WCMSZgX77pwjEwX75jmN07cfEIu72JJMVHITS+g
tbsYadX2QYtvh0WBbhUejJMQjw0IW47UAN5ygwFut4Ly6n2z+Jw6eqgqIcxWM+ZWOCwOYII40ffr
leYA4vUUX/VCn997N1bThkU0wt+eOKA8ieSlWGMi0K1rPUv1YfdfYzzE69UgBZxijHGUfm/ixeoR
tJY9ZyFB2jz/m6nqHMM3SV61XV9HjUxyP9HEP15NSwaOmaHHRqakppLL1HMIyQAjl2ezI9g3NX5B
c4HkuZK8yhMFgtfkjyyaSdFzPfaaBvx8gXOaN6ZgDWmAWxngSpEgOAHtrLmLL4RhLdNAcfX8ejZD
2Mak0INVDN0e/aFhH1P0LF+PJ31A4c9sH8idXOnT6l/Vnrep5nWaGlaWiO0VRSYbIgfjouml9sjX
YmwEe4kQDTgYtIHwj99+2aVK+5mzntpD+RM0UTQk4usSwdEt7iXmIuByFfCvgs6eZT/Y3w6btPYf
ZDy8D/6EC53MLlxWDfvGZbRssvs9GogjtKs04Aye6X+l2Dx4XKxdcKmk8VcadsGfUqrQKxT1CGgR
6ndkcW9tTyLEhVr8LB4yGbohDR7DC6xO30mnCunb4e6uD/GuPlzH5rKViXDZuN7hv/huzrEIE09c
MTss+HHvOyF5sjpQIlcLg7b//mSr5mKInjf4g66IIsmk6cG7SzbExnlLVU+cj3S7zeWP1LEi/sh8
xQDwFox5GcAi5km6O9ySNpc7BvtX/A7B9rcy64Q8x58Fv+7Q6vLM/u92vYodQ5c0jz5KoCrOrlXe
aacqLPzl7Q5sV3PX/E8w0dBRS2ww8nj3gE4JyPOVLZxc0iUYJjIvomr33bp6Ehg7HcJOoepBwfu+
IAuf7M4NMPg/dfuf0HmlWVlxeutRONdhQMu/eHTe2GgrGRn8SlrEhTyPQpuSLZ4jJaomHJNo5qEd
+ZvOoIY1KTYUtcGxMNO9fJaQJV8b523CqwCai7pEopfBZkeP8YV7gSHJPqWdleEUEvoALSABuTAn
HCZHE+yxNZYk/iF4y0n6kiv22NvA3UDrDWK0xvAGlDknrDjVFE4wqtSxmFyZaXQv86CNt/2Stx6l
hj/pTVrVNC/eRdiSLzgcezaHsDyquoozx4tJOYIPmHP+wHgRxXQmhIBf1cZahptSiDUwU3BtQTfK
G/Iss740exd8/od0FUQzjWF6NICHl6xSeNVy5DtfF3A1gabMKw8C5tuiNhECPDGNko9kXiwAGWR5
YzwrI0hYo697UAoXQxIQwv00zws/nMFjPavBnO4YW4QgeA+KiPutOqmQdwQnq28z9i8GnCwT4BDU
G4XQss2mMlPnydEfjPL7cZiNbX3mj8LiAA3hvxZmdlEsBFC+zS0SYAUxuDj1rAwhLdUFuDAsXazj
4WN/BusbhvDB6JXq9VrFN2unWTC3QM5ZgZeY23AuQUJiv6Bwu/N3zDbQbnVWUyZnFW0Dwk0ehlqm
oXsMdOxPcX4i3KTgDf3366liLXdJtsQUD3HnsZHWjFS5HuAazsUGxd+esShDjPQ4rq7Bv1fHrzMw
RGoe/HnMoZvNXTuenuKGm4bMSN8qDYwsfnIe9BI0wWvmjGVlQ6O+/d6yz3oMqPvHLp22XL9e7Es2
u7gHAljUhoPDJvqArrVgJCEG/LDWfzXLgtCAl565P+luZjTwcDtfK0IEz/plHbQHfbeJqeSJERHl
9F3AUIGm/CZ3eObwWaQI3bcFQYEzy44ceAQpKnn6GznvFkR3yOTDytiRE2UsdlPkmsuXKjOU4kmX
v6IZs3W1WxVPVZKXt6Fk3fHgElqXaFuWsWhfRi8hdXAVx0Kh4lOYQ4PTj2iKh7yQ1dlUySqYfchJ
z4TXvCkVFTNaewqTuEY9u6fWk6HRqJ5r5oPFfuH9WYqjnCPnpUsuajrrmBAvNLleJPTQDdifMr+T
V5W21vRwMJhv4W2cyqFNg1Qf4GNSlj18M8PbyHO/u7vS4Hq++WDUoMj4kFFmLzo4liC8U/QCVJXx
xEPflrr24RdSpBnkz14bO5pRL7CBcy0PwGym4oPONLIrybLpUe0v/iLUuvXnGka/uJxapbZbunAg
FxnxF7OI7CV8u4V75N6aD0SffZT1zU4SbQrIx9mqHCx28aO8toFRWWnbuQ6izCtoWDBLpNnbq1Cy
4d7GwrFnRwcaazkkFGdT/LhO6ytZfhH0XRQ+J6iwFoBJLwciawa0reqYr0V6X0cia36Oruwpg64a
5sjWprBiDVFCrzQScgi3v2jSHPOUIZF3l4bpjLzdNOanwMPEBCutbc57trBg66BotJJEYtzU+WPC
oNH3UhTry9o3rKTF21EdY00lDzf0j8qEw+5N/Mfm4cpPSJwwDF6cbB5OkDwx07sPig1kYSXpF+Uw
MMhLMXKASYK1d5fTy3hO3aoRlRUF//HvHxUkTYag4H/PjvLOJMsY8Ukxt2XJgoCWBNjMynx9BWze
7oht3kDZuZUJtgAGXzOK0SRffzFajrHyrQw5voDYeMsK4lQkgdf6Ms2ZdtRjZUYc0rPFfEypbb5S
fD/ur0j2yJCp3RcxIszTtophoG2AFGjlK/qavC9TB+AnnJl924BgnAWN5DBFvZ/KLQpwBz/+9tS0
VKeXLUozhfBjnYqFvChoS+FO8SN2V/j6pM0oU444igFGqwKJ+BN9UMnlsV/9zgavdD9WDA0Fvm0t
vc3/giXvndXe/9/SGs44dkQHDOmWlv21cGvpQ1DTy3rwZl1TFQn5J4V6S+WEdFN1bCommR0LOXT6
RUgHCCURVPJxZIE+NQ5U7Lfvc0MQT1U+EFjHCKDtZL3KbuRv5pmZjM6Rm2gTDJsySfnXInn7+T6D
cxWFSYmn61668QYc0pQBu/TnVjHVOQkxG0vEoQK0Mhjbqs5ZRfpPiFQocL9S6JbLjId6zcFgW2v9
jN6mhA0Z7/n8jscQRi5fN6hQ2xOlbtvsU6+6kDyzxrNwugfzHO70l0ovLnJkKDvibW08kQ24oCM4
g5fBYJ6RbSfIkkgd3VaGH4yDcQhXNjUrxsPfTqm5ZmkjLowsjth1WlifcLuqJjfqNUqJJxfELp29
BW5gGCzJN45rY1CVXfmEuZzaHMmgglUihlLk8k1GKJC5kJC7j1J/ASCcvHkbGbSmxBzKFiyOYFIb
CrXNGZIpLMItgroQnAw0HHb1NTSMMy2yNcXEXc1fZtrfnWTJymSmwfogL4q5IghSTGC7vsBg6Xtg
O3RQYNp450xPt+OjqEiSdBTLtvbZPCv2yQSf2dBeUuuud5EK4/go9SGV3R03+CZaIuBaBLGyPjZQ
IjR6subJBoeD0H8keArH3aPxqUH3y57MoXboJ4jSWRqYBJa9kZQ2UZIiAaqoXo/SCLQF2jCiWTjx
qDhQBBHW2ZUmAJ9tcdIafBKISd6Ra3s2UmIOIlYlNKsLMEE9avZDLT3iatpk+h9l0omIVC3csJaK
z9z6dur9ky82AxjndqktKer7LMR1Qdjn1yQuVJsik1//j3ZUwNmHYHgBW2tMBDuHjpnaS5LrdFBe
NuXO0amD3goVjT2+A7bEZ+Hv0biGmt0X9Uffx3SYFps4mthSWX2K+WoCQIOk+gGlmELfxslSfIVU
Ck1D6QlMeJ4IxJ3PMZPC8PoFLtlbwHeH/Yr6+bHzf70zOkAZoA6B7/TBJxooz4lwYDmNT1PR0/PV
Ok7XdHAKcbkOwifFZUQoHZVaXngWk7t/zHLv06+iRW+8yzSMI7AT8DnDqQguKFTHnBx6593S4wQs
cZcTE0dz41BAKxwL0+mtBcx9/MD3QQG8A7EE4+M88xaZf/fP3fY5Ocpp9Q2WJ1txe03HU6vqm6ah
4J6jx3IWBXuCtFwAIYbfIZGARKyZOMHGqF0TJ4JGcgrREdnMoph5sIu4PGi0QLqoUb6DqwUir+Jq
bTRnwzJPcl/Lv1cKRuJKXnIKd6IguFe4ddFVI/W2sHz5TMrgkQVOMDnHmr4JWjplOthAz/dYClo1
gdJjV9LjOMDxrPj5timJZMbqEovyq76G3cJXSug20uFnNB7MsnlN+jvIMNaRhWa0Adaw4gl/ZMgZ
Cki3vNW37vTxxjOxD1NjfnQqJqE9Cvz4YaWvdtF9miHcxa9h5/CWxdJbryldAWpgzWE74a7eBAQI
6CIXOb+ib2UYy2tW86WRMKmX+bY1HBKCU2s7r1SbksxjAuWOXdsjB+LAGMd6zqyjt52ne3gL+IWj
Kpi4L8wpbdhCzHSm2LgzZ4CsakZw8MR2YbDXf5CtnAqck1IFMC/KjAigRqPFH4SJtKArlWp/mhDv
tZLi+Y97GZYjyhy+SYNmt7Ypv/WLbxN6TUfLNm9SD/3BfJMmN/OPg4NPfAdmiVszQXW9YRF7aMUe
Cw/Qs1BMz60u0jD64Qf4Jz9cxM4XZ0szNGLSdi0HcOk144FJo5za4YZs+8g6G5QFfhuR6oIZNrYZ
Fk8RCt+5Tf9TxauJON+guB39URp4gTFizUiXvk+RV909FOhaMStGMzuhnJe5SAuwN4YpKR202tUc
HYHLQCKIm1keWDS66Q0mquAHctDiOK9nlz7ff4uhXpbaRLhBXi3LxX7ga+bPOXzTKxuCarrUj0a8
wz8umTl/JjZ/joaCNUeK52c3kRj4SXoHv3X25EI4jRdqc8ZvfhzHf4S67zjurspkoby2JNhVoREa
FYi0YjcfdMTfBeNs/DiJHar8DkZgo9N5jfslvbICyXm5fBEOKgPRv+9ND7HqkUZ4tzmojDI1o9CU
frDuQ74mEzqiZHRm34ut4qmTc0xN6KUNhNkGrc89tzxScegYnKh//3KLbug2/pXgqv8dB1gOuDPj
qwre8dEd/OFXkbTcMmVnm4vVCWXYUSRXFgnAB4rcgRhMwYKC9+e5oneQ5ro7YLaWGd0NZjQGbMht
q5/CbAIny0XEz1/B1I6S21yqf8lC8FWSP62m2l8SNEK/b8HC45cETyBW0zT4ZrmhBBEZWBQFkVc/
HGzmeCnXp/6UkX3S9QYu4DhJYSDDWDzDR/bbHUHShj+0MT/bYYakyLT6tJI4cOduNLYm/DIGZsTx
HsXY09m6CQHeYnY0tyYaXa/3tHsRmB4Ic5Qoh7rO/6ULeaoHPvMaeOD9GUAPJIp5X7C3vOXNl+02
Y3Yjm9IdY/yHEg55eJVMXuOmREmKNReN+eL+8PqmVLZ4JyHk/+04N/7zCISNEXcPCZC2BQG/oc/b
Q0zInHD5ITLefw+lzrXV6SF2tO5WLmZwt2T63KeyQwCvp+0BNPJzQwNBLTFk4xvhKM5dxrjRrn9z
syasgDwWDMbXFP1EbVCcq72gRyjhMajYN2/hTlX71HAzhNBMyVF8+eTJx/kytClsaXKnelBlw5Nw
HP+RVRd9gLkNQEw2xyo/QU1nE4rEeDCi7WH9Q6dxU1HG+0CaUBX0SDXir+Qi5z3CcwyBTNdlEKdu
RZrIw2ZUKsDeIfJuVl73RQlTnnVjr3qCnUcg44Ficayk5en44nm95F8wgkv6etBHITVmE6USilxY
dsw7AnodJWFL5ZtURk+CS9ebHvTOUpXG1b5TnnpQ5V0nouMSZ9r6TFlQjJ7+79pqHUkn9QgEA4XB
8DWEB2K2U3M93Uri8PVWCZXP7LKb+OGM+hyaJFytKrhu0m7m5EDaXYq8cjZZisEKZJC1jBrnsM0G
I/FQzVcXoW3ObPp92jYE7UI6m5DYifyO9R2VZWeTJLxXzfuRetDPVjhtg7eqptQ6K9Nwn3NniqaX
ED0CcKt56A6iiwFCPIn0y2jM0UOFio2/9zMTyun+Og9ByXu7uhN7DpqhZjZ3SHqmq1Y3D3G2v4/f
OETUSuirmTb9yWSFnx9BDjjCX5aEoOF4og5GEkP19I4GoQPZ/nOa6KTWn476M4sHbwXSeNO4Qta1
4DpA0FXOjQ369C6hORlEKsfDWZgQLivbuiSaWDRSNJoPCzLBRfXsDEg7UWKc7enEiCoVjVFmdf3r
FnIDUtsaAbCT8LEbec0xrL7DNYDC1/WwjsfxKNnJ5184nSTKKbXeVG/lahP7DyJag3s13DlWAwLu
jWjqMYsaBN1qtdK4eD2wkYfIsNUDEfyw1pOvVw1RjQnFwRPcTIH4L117wbeDPpDER6CHez+ZP/9R
+C2WWk3AksdUYdorogh7TC0gKN5LMh/3yda841eHTLsSXfeOxKeegYvzQ3I2IEYjZ0WSTKfFd0kR
kihlr1L9Je3mGxZtDy5ENLFFPojuS8jQi4FpGfnkXn3J8Uk8YMCRhU4aZCC4KQcHjmAA5g71beei
Zn18Wx3y8w1m7BLmINk0JfYyppzAdWz/my0IBwCx3EnB2qVWzKZVdjrsuDaM6+tHsfl59Vby2jjG
BCbD8nN6YEctemZKhWXTtD9n9HRArfcwggQCorBnxeOkjNv08fOoWc0MnnPCyMjIADv13SLC5qUr
Bp/F5KUpbSWygZPGmAA7wFbjVs57G6dPQqLSje8RRrnPcQtm7BBohB8FGrdOk5XrsrJYPU0eS4Bi
98aBF95FtO+kTYKQ67SOInMN5vE4a/sFvtg4UJ77fQ4WMyUJtmx9bnrFe2f3+PJpMsZL94/camo+
hqpgikDBPgylMSLUY2Xl4lK3m3GeItXr4gHW2RRhLlvnUPi/ee5kKrVcSWlcxe90mWN/OiD5/sEw
BOxFxlpgDIx1VJQ21Nk2XSCxBqh+Oaowb9GkytGhvuGEYUz+dcQskd6MDF21VYGKoYKWchCAwgUd
6pKO7oJ8ekl46SkmPsxY26GR8COw7aDXrCEYQqKXvXsZVircNAlJ6HKtdU1Hi0VEe8NlZgNwIYi4
bFHP7P2VpoPenlX+8JX3yg436mB/rXwWUH+wweVIYaJKBxCc5ZTMvMmSZqYBaeAv9rifhcIlyAP/
u5s3f8MSvygufZuB/RhoNiPrvX4LnATNWVB1wT4wPTUgbKYqdVrBtQKlP6iJBM9nGWlKkBqRuV5F
sqvu2xuiD/ViQjMwvEeCyO3P3Aqbb/ECtWQOttq5zOm3sQJr+EaY5i4bMHWw2pIO6ykDw+FPcc48
NV3ys+9Dl5Vxut4tr891bUiDUuWGbhM9oi433FnFMgl0DryHzntcy+Ky6GgBw5e+Dn+JRr62eKrw
njhSaETvwhqQnjwA2LKeJxApd6far4jBTUe90gzCkop8Hj7lAXQ4MjWHy3cOZrDLJdJ1yX2smjyd
7SjBKAVbOwjbmCZx8kFb+JdDJBwwDWIW/Xl2SRX1Yhv4cZ6jBUlyAmq6c+oqSVKPGJGeHFfgwHWR
3TvD3nqKtP70KYPBA6A6Sa9pm0z1k3KAX2Ze5LDt33g1Tw+puWyNBh9haVDG33dAUZWFfNohjVJn
9jC+scmzpcYDN14fVnJaAzXcbxA7/Qb5zvJLAuhjuyk7qPzR/TWLT40AhW2V29v1aWDWFG37RrP2
TLL9uk78OAbWJDq87KVbr5g72j0TuHnLMR0xjMNtQTHTVjES4JwA9TDXcQ7mcszJtPu3hUSPSZsa
5oHlwDeORGjMCCIqBko61IPTEgviak1c/d3rlBda9izxErQDXvMZl9bURIgnKPrWKSuWC95+pr5R
6WVpVN82TAxAVnvoMXf+DoUhUfNl9+3iq1X7JEJIlLXIz6ocTbtBmGCUNs0Aw1zfyTN5BVHEKxYw
8z2y1APRWMLXYbBJx1k5yG1maMjhp6MgZ1Y/XUcxeWt+Dz3xW+NII+hMctnJmoEgnPNzJJLCwmoe
JcNwN5WaNfk7oh46v8KrcKF+7Ohqmwl+CQsOeLNk9B94oRvABwpbNsegr4qEUrBLYFOJVaG6jSIx
t1qrA7tppSDr4jgSizoBO2idmnMY0pF0kKeurhWaW5hbXWeVnq/SAhljsjJvUbM4oI5uZ1eMyCcC
qAdOUQdNYEh1zidKEcVcZpu+W9TEi8T17CYyPh2ENs8giP6xNe3qzGlprZGZtsMnc0fzjJWf8EB8
gdFpdFQWc5hx+wKBUo3MMSKZqN3LY1RzWfE8xBXDXwsGz4VN9tHJ5zLzXkqOHxxKA1Tas5bc/SUZ
D0zYSrDqdd3LXiLnlPqf1BmZxhQAycCxs5sw2u6pVx//TPIPQiCi9wDIww7y0SmU38KNCBsN2a6S
4Pw4FdZjfSgNybhI774QtgbMkBSAzEyXq74A66KpOgllnY7R7WMlAgRUQNKmXgf8jK9smEX+aPN/
R3K4pZoGpG67elXhDCwek0ZhxHQCqv1T22rXNeezvUXmcoOVt8F5V7LX7rhLq5qUIdJfHxm+bNhe
IbqA/kr4w2cO+d+lG5YJc1YxCwmadWthFfvbuxMRKCwf0FSuNFJm49/zI3Wm3a9fx+XY9qUuZSlT
XXMIlSaVh0aSalAmkXBc8Nd5GQhVE0t8Zj60XeVWFjqrfXnZSInI4wlDGQiQUjwW1UKYhVEk+i0D
bH/aPBJvUPW3UDo9Ja3SS0aSgqPALZ04w/cwITMb9L8EaL9qNNR0Gze7JzAYRMLW8PyOtkP/pz2g
Fun9VIH8F3H/LhV/a9fpJSn8aTR9PdQgv0zFaOS41JwQBOrgCxD6WUt2iAZj/8RqEsQ/ZrHwt0Hr
RKvj+Ts6/6l4ieV9+MmKxPx6qsUhmu1HqeehxrfZiEcW+IDAgh00e1t8urLV++DTR3NmPuxg2mEq
HeKl863G4X1+IUMPDU+dLD2yX8RJ89/0Gi4qrP8rD8Q0R/GDzIt0S0zONfjHByDGQWTBd74RdLMd
XLTll57DCyx3fy1JFehUZ8S/0q56q427GmGPkdV4xmTApYAKlgW1TjSpnuUAOcx/Yr61u7uadeq2
ZuSU0umIDGDbFDH9wcPg0rZbN9eEDxNZcjMPY9k5dHtWGN9zUlhmHXrzJSG7np1ra7CpXvHZ4Z8H
7RA8sWfvEYYCSCPMZ3JArDYKL0Ao+eCx/4t2FfPX3u9QrX7X40iMNzSULjKaarRlYV3qSlo1cXB6
/9CuPlv03AF0sdL+aGCbhS2f4IzRlNc/aECj7qDrXltu2x870qwrUikGXAujENmW9e2KsNIWyYeM
IjZ2AUpHhBd3S/bUGZoS8cCfapAUjE9d8RtiAfzZ7Sv5iyUWmbXXMuCJqtpCWieycJ8OQrRr8hOb
j+qYOVeleP06hL12PUiANNFiyC9m0l/b0QJM3Z1MCZJKyIitthv4SAqWHxL9TSC+LSZcS1KrNbaW
DpVmYAcwIkyFqXawPTfluiQ7+VgNJB7f0TPg3uKNMWEupGSStBKfc6oudGX8m4wEd9hCI8L0zkNW
No3o9DKSzvfFj7c4GQE4aweypSpH16yx8QlCNQwjepGxXAi5pUjChI9wj7YJi57s3LyQ0TArvxmd
vsrACWM3UHBCy5jMjagSwXrPz58XDfd6zXplodMu6u6J9n1CEiK17fAUrYiHjx1OgDADjJYgSoGZ
43UN6SRP1viW5fpoQRaWIkzvziVAT7cECBpu1ccslVGr459dKb1wLQvQ9e2BQ+2RVYXXiGgGNi5b
yZ6uH5kjAXcVcbIjJ90jYKB4ZQ+AaYpOvvgNp5P6HFoxLBHyTHCb2wH1XL7GbdvnXsclhUvus6r8
e7xzfRZinlkIZannsSYoJf3kbJFarWfkVqICcu8imB/HoBJhr9h3PBlV/ecL6HFeIJp9TgY4VeUp
ZQlc9l9krRYc1YR5F6FFGS82HAYpyuiWatJpymkdVtVqXWsnislclprt7ObZOPmequu6fUR18Ep1
AXH/j9RqPxhHXXi1OVLub+//UTGbhni51PiD/qSd6naEOJWekbHp4X+240GOrqRp1pCE2bT0iEEO
jxfQbX+JYB45KAFG7llk65IkP1aLWE3jrIKUpPVYf8e/Z0OdXmE40cW785pcfQVT1nicD5fD1MnI
xysbDw+903lZVCV3SZxxjPlrQYBVghMOiaUBgoEoiQPRBxBI2g24rrdi1cOyGnb81USpw5+gQthw
VDMrvj8ft9Oi28uInmOPf4qoVzX7AAdW8IddvzFC+WInbRLTE4XXIU89xox68NHN9OwRdMG02D3U
Fmr6BQhItTWHWpWGI9gAC5HhGqgCZN3+grYIC3k5KHTRytJ/W6EG/hFli4qNH1L1mhQ/GkLX94DD
RAcZQXHxIvV0TRcKH+jsJbtn2G4QbhHii+R+kyvOePbOFIBXDDQbgkVbH8XasbIL/KkyqPlXESZX
1tNsxRpQb1uTmfGetVlFzkoax6eSs8Abv/ewxuS+2KQbCfhBRKM8+ABzQ4SV77FWUG4Q5G8lwXS4
S/5QhAI8yA5toU4A9T3Co6IrLlJysilGkwv7ikmVIgKe6rqPfXWJ12aHSV6HkKTFOkyx9GHsnuqg
9zB+scGRlRq/x3yRh5uxeAVMtkqd9/LVpEVjTnn7LcB1aYdQfEtOOF2B/GaIk9uipKhUniLmbfh3
ADNi7LAd2Arhu091Gq6YZpnRNZst7SOXpDQfwmpD9fT3RffUFzkRMyOXl/lH1uBtljNieL7l78Fy
Q2H/t/vTUhsEjxnXJEFr071o877dxzy1UXTTpnbhi+fyOXHLETrzy9dQnxFJVr6NtSag1Mf/9Wa5
rI6+N50zTdqB5f0YotXmfwxKLOpvTnkkupVNG1b53NK1/SEWh1BggG94VVKQoVwIgbollpnd0S/A
EkDx98fkzL6Aa/gSMXxfEDFzJuj6ChzNwy1AN5QkYl/9MKQZbkB8IiqvCw4e6TNOjcrACv+Rnz5y
wz7ZnhWQQ31I9YkB1bOiOH/6gKSKp9a7aQqnLvnBuJCd2tUJkP+qHxGtm3Wkb7PUriHMvKa8akNq
/Z2eTlY6XBXmlq34ueRumq/8bZ3tae/M5CNN5MOK6whEyNMGGtl+qcIhvDzV316GD8svrgOybCBS
/pP/H8QiiXL0LDexNYWzK99BESkU59qd+B0ObhNaUNQqs+4cfkfuo0QdOpZ4w3e05eumxSrkwqg5
brAUa4eX3mUfe++Cuv7wnv3jqrlRXY8rmosGQ5eg1454U7ko4yK2YuLoxHUn6Kikvc5XUN63Cdww
sKezVUpDWp89j/pjqDU/d8e7XT9sEuRiquxgLxgIjRNG5xBlnlsXF6WwFq9RRhXqM16wlixtYTCN
/IbTQoTieQu+2eL4BQfD4AJJDfPMu4zeJZkgqcTYcp4ueeTKIRlSI9nBkYo9HtAhQsSruM+r8BPo
nltDrl5qoKj49TjXbYH8DKT4IfG839LcVZExGNjDCuODUx2KL5xFashhbqy4xSd6zGBv8ZCocudP
5Ck8Uj0OdVH1SgxWRQSKzmP94LWwv+cClmG71wL9Kq8r2qU/J+EM2bs18cjsIcWnYKFgzmr8Xo2R
Wxm8Or46n8ooyrXp8KZM7oDNtMCnhwBfA7Ajq0NEGD+I8QJEWQ/Gy1Mr1t2dE91WfWeIvwArRUdy
1qIETSMz2hWYYQHdpFZIKL9gjEFbSu7y+slmw2DDRnLyaGPlapygW4fxfuuDCbb7WF0Zi63JDyfI
/xr00edW9BjQzottTUmNBAaCk8ogocyKaKvG+yqDJV7wmGkb8+oLkProqOazkkLgbrCGUA+iX3d5
7yf2zjPiSKwECbEaDkHdjXG13PmAvdNvzE8Xz7+JKgwzEK8z2k5eMtwHx69iQAbECk5p+uSmurkg
q8OgeV6AZc2lw4r0OMCgga221KPBoCrDWm1iKZ6MunWFZKfjLRYy4Cwcg9mIVz/p9Oc1cXzpBeE8
ui3TCfI4kj45M5f/mgZtlbJQ6SOza1fnCC/Ppz2varkIUkvfgJPYK9echAmlljNEOD4va6p+uEC+
r4wQ+eEAb5WAJY8ZA8dEPGC6Ln8CFyWzL0/lalfuSJMhHWSEefVMlbB4nX4khKv4DA5J7+PShibJ
kof0KuytEJvXoIzcAz5sWllIshLDTbL1ZJMgiOZRl5Z/dvv3aVyGUucCksZxUSnlj/bwB+VP2/hS
KsG1iakzenIImVeBgxtQM4nB0MMALPl8UXdCf6O/buIXYtZSmGXcdzgly8brkxadGbjaFKNkmD4O
x9omZuJ5PMzWyd10awkJt6RfjkCz5LgsfIX+dXcXBVAFpHa0V31mGl4q4cw+1kYAgA3m5wEF4i75
ftipvyqMCX2Bv1wLuzdItyZJGtCxMxPt2JC1bMeQAmTDqGMXHcYLOi/jx1/OMVzAQKFr1K+P62t3
zkETOeRnUW4tTGxblzyp/TcYWIPnATbRHZgGhWd9UTiEoXDYukbbISfIMaH0KK4agoN6vTKS0jFS
m58BqFLbkN/j6nkCtn0BQ4RymIByWGfkR2RKHsZPpnde3leMuqVLGkUnKM8Ae8sA5qzKmKKa9BWe
XG1MabrlqhmuflvBB7dlDLaxtvEkljWGFp7QUXFGYiQWuzu4Wg67JxBZFpA5vVbrptiBlQtkIxVt
brBojyV/RYxUK6hJhXuIVJKi6FGwuPQZCa51CqXCwWOGOLdLSUJCOFPE1e5s1+Drm+i3S96uaUWX
xTcKRPKZNtQxe14MqaHCSeWvzj9ywnc+vaczDhyafpS2U3AjaTfveRxzfNvxcZlpusz4trpz7coH
9mR3Y7Y9F5WsCP6/DB5Ib8HrRPNod8myqwRgQfSiQ4j7p37FKYPWoOy8a7AgPCFi5A7f581luTBb
exU4renX99aZ0oNpSu7EixjTpClWn9rT8isBA5EwLjrpGx7AEYjcKp7SFJUrSXAwUWk7yXL5SDTm
o2ZWqCNV40b6/+WgAeun9Oqd9efPdc40JmOpCZaTuyZJAPwrFn2emWY0t72UvQB4Ls0oLVdSkAmq
LZQc1HezwNJyAdQ+3bUb+kCWk1CbcGU9aE8zAvjJ/8G7tFoamEXNZ+FxOuCF4DgMBiACB2SK7lNy
WXLFwhyFjZB51pGVInCfEgh0z0pJaxjRY/ENXjodUwnseU37NDgYgPIYg+MpO/oCYIXy3+eOTDuh
CmQ3POOY/Yc8X7hxQ9c5HFWUBTChcGi+F6YNn7zomLG0tx/oFQ5t/A+dMz9bSZJ3fpBTGVSiq18E
rLmoztxQzD96T9F4PS8FiKwp783wrh3Bhvv6zOY6T14UH/Lt4VvGWSx1YWDmrHdnBtBCBec49g7x
YpNLIun+0gsuVwyXUnSl2PsBlg4zmxKki9KsHaN4Uvj5DP36TT1vyj3JFtEf7tpEwl8yY8AcN5bi
Yzi1ccOYTDE0s9oxfv578xxcAoewxMkQJSZV6feEZK2/kLqGx6ZRFXza9YPKWrBwvDAK08FAxM91
AbwE3O+Lp9bGuANoA76co05ka7QeXmiU+8eNgY+peKZqrESBvOKGpXXFugWxae6467LwpML1c8YE
9KSq1iYezj3zZ8wG+Uu0d37rQdUua3yuXtb1W82ywMXbmEwl0M7OZTfSxBfRgb5OCUC5HhSltxVl
sZABpO9DdPzVJXZcDjbNTvdVD/29v4Jj4tom6VkZiWBbUFxcMSM9tjFWIOd4UzLv8UPmciGBPztZ
SIUz3+FoqRRNTiYP8gaVZJcNQzVpLd25bWt2LTAXIkz8T4+/qvxyBUKA5hllXIraDFz+KJuulPOl
yuxQCX9KJ3pyLBTnq/1woPYFjNDkdcIkorHfEFL1/bWARlsLn34QNq/ebuFQx6VVxBgD8BGVwJ4Y
Qe/yDppDDhQR9qJSptzE+KaIOVvulawnY5lNCI9Qp0/fvMXPBJ4D0smzonPvFdTgEgG+lMl3wz3A
41hW+GbETh4ubepCZuWSM4gM3K83w03yM5m09XurY+PSpzVSRrm7y2l/8R0bfza7GIzj0DHGEuWh
Maz1WLCjSOhostwExtP0QjYD4CTl5Ygcf6R44aq45rBYpVVypaG1OU5YF/exyNdkWLJy95lTFYxJ
WDePop+JrsW5W5pi8AVD4X87RGG/OAgyVBEtvZySJRQ3BFuR0Yd8Cm54SBDe6EXg1cpW82NhtG9s
NQBNXzyE8KoeyZpPbULw0NMtpaCXGTbeAr+KgnW2FYoieBpY0JJOntctdMY7gLohg2aiWWOxwdGV
ufEk8UQMYTOcIE+eNiQk6Y1I5Dtfmq5DJ5dJU8pD8nZccQTqWNQbGabkEk2Rt60jQKaFuDFqk5Gt
uJ1qh+/mWuSzEJl2SPmE3zwKeapgUG8zPwhmW4yo4CH1KtAOvpmvvEg3eZewgF+Bk+C6PkKl/Zxw
m70VM3Yb03gieMkH/KAD126npNnMRqnQXj9QmIMiWUn7NEePcKLbE/91w0AOKJQ6R3qMh5NI2db6
xCuy4mnh4AxCm6l/RZobdPwZu9DKX5J4Pti9J3oMYNhLHYAWAXZovO4zlbmYU3pQqZpZ+sTT383e
TXqmAqU9q8wscMlPyZMI3P3mwDIgTk3QPSilaOncsKbIv44LQAIPuodV6xztSbKU6lHQdDPT/JQb
vP3HU8MxIlm+aKpsJz15j4oRgu4kuBMiQsm7tJttggr0tEEn7U9jRbRt5u+7eu2FXSL74H8Zrj+a
4OrxUaWRhc/+w0bH2xmjStB7kN77c5VPaw2qWaOfBQ+kCE8JZQfaew0wzLeOyZ8u3YEPtasZZkd8
+dPzciL3MMetbOcWOFixbxgK4jxqYqHY8Qg/j/pABm3wNoY/Ef6Ul+hupSKFq1PXFPN7gGizg1wD
kxsON0IcoX+eIx00WU/nKBSQ3z/OsoE2oV5+wW1DmpuTNXvUnq289S3GVqo+FQ1kwJiMaBAsZShF
G9wgkvBZc9qgu6E1s86GodHQ+J5Cbtf7XFbTeDIA6EWhLiDrbdf4CYlxl0UqBFgQ6Q7Mwyoe34zK
cOSaAiDZyRhYs8POJT566NbS6dToJrUcd0kt+iInCowmStV3gOgpI6K0CuRU0JHI1CE/tpr2fDLY
rOIpV5ork+dsvsV4UAaDHUGRpAyb7pEMNaGd/DNkUaSKiiA95kVCbSbt7dgcJK34iWKqAEUijdi4
yIvJzVpqt9+FozQzHFhFeEu1ZqD9eQik62HORFbnJcCahhaY3mhw2qSVoP1URGjNh7xvYzJDfjwh
IOd43xvXOsGtTPkI9/iNICX1guyctHatobM9wzSZAPwUoOAp4B6OAs29nV/f+CQiIn6pmRAjrr0F
ATPXDCVkIEjYapR3OssHdkEu13YCbpS5dcdnVvki5l3GtztebNrrRSd5sIiYtKedtVfhQucBYcLX
oLIg+dRLFAiibanRfOAS7WJ43rYtdRmY+HFsy75HP21vzZD6afrFt7dNVHF2jXod/mF7qbRpsjR2
KS0p6BXkCNhuM8o3uGadXwKzVBCUDnMRFcqTQbtTMVSBnw1uFgYXachz3peIy0p+HOcbEyyrJIMe
iGWmjX10TuuEPNimAeS2oOSsTaZFso0Tzh+uiOfwGZmsrLYHaRYYmsWVVh/jkMqKpYFVuFkpqPkg
Rm+MHN1r/SquQh/VE+I1q5WlK8ownUPpQCa8QeLesggX3giVSCkNHWo3N4kx6/jugL/P9Y9D/k2M
OR/UJgNDoIfWNWaptyKrTQvGdZWd4S23U7dZ8u8P4M9ibgafz/H5mTJo3WcPCGAYp2ZfJA700MKS
l3H1qBxAkKkOw6JoeJnGw80YMeNWuAOFXn5FW/6xReMNBlxv3O4u71FUofyzKPQoPpRQcyY85T3n
Ye2bwg41PKVoAWl0uG8VOhbxMPnwDR3gnK9QdyIe+8BR9axq1epEe5q6oH/SPzpmzYrJuF/YRqga
wmHLrby05rQvGUyLsMEIgq4fDvQq+epvxV6Lw08HtXQXClHgGpyaEfgJ7MyTbtxKk/8ySQolh8wj
Fc+K+ReWgLFiMmyQhAHFy0tvwrREsz1KzRM6yXDYHgwiMx/RMPBNkvN6szxzr+DwGbYXiEU7Eiqh
0JkldOmyH/Vcr+GB/9LCDgRmhFryJtEz3a8juqMSNEjmeteeSr6kSTgoIFWSsfMQ5B0Ta55Y/0xB
bBa4NhyKE0yvZnZG5nkWkZv++4UEvM42+yDvpCfzQizF8Mvcs1JX9dkKxk0vgNB/pysAp0Qxc0xh
6uMpZ2EfqlIiBWvCloYBllbPaCbhR2qQ95wSxiEsKdxMk+OnDd/ovha2LULmx2Vi6YRIBaK+fgh5
zwHNbf7aR2jWGQ0c0T4t1ocqIMGdtjhhia0nraoqKDz8nJcP9HmTUhs9Dz4eUDfx/eFtuu5RMym3
qLq30xX34XkY5JJUUHKRnK3+5SQeYZ7uL0WHkxKeU4wQprrEjFKy3WNxgtkcUdefMJLKDkEfrD+Z
4LBqfWouSACJSD6O4v43fphSLUE0Zsc8QmLeIBFnU2B5fn8LAmDdjg2/UxpUtudBQaffoO7IvHgx
xnV7DPR3KqYW2kTT442JQHqk0pzCeBwSDNGjUh8GtigYxrhY4JyDj/+zRCpjnrBfZxuz6U7SO5EP
Qdmc50n0bp2mUBU4VVVCbVFa98OcbSLoZ4AFa/YrLaj7v/M4m+TFFLo5AzinqJtyMzshkVMlVqxL
yZO+h9rjiz1EVHO1xFlpqh2/8gnhB92lBu7qW319qPu4QUKpxQQdxLOjdELC9AF1s5itG2FHKxGZ
hbyKXrLw8Jm/x2N7ujlz7NUqRbbA3YKiPi6xoEBO5e52M5K7dgT+BA96ZTgBYBVHZ65Kw37VkPGY
aCZ8QUJEg1QRgqdccvyP8q6HTK6NvNh/VyKILWHU/PZd0OL1ozYB6SgUOQ735reN/KgOxlpxW5fd
sudx/ZS+4nndkb6d9mQk76XIRw8QC7SLtIQeXm40y779MZmfPs3JtacMZrSNxzrpwJIRAiYrbMLp
rNoCdqdDVyievMGhba/t9j+FK2EgzYreCLB/gjHDPvrd4q99fzzXKAKnZDMUokAhnkX1/GOYVO3a
7vTqeUXBTmduLdPHqSZXQ0B5VZfpcZM9y3Awb0UDvARxQysEVW6Wq80YRGtxH2f+ulAJ+l0Ms+zQ
wOuFzrt4wZrYOtTpC1Lf5T7k9/Vps0r8lcmW8+ivVfZhZuOhRUPQYO3/bjSoHDOVLK2vVz74Hzzm
wwHpoiCJCZZC/2yuJvyPFXTjKH5gim0bkUdihGVmGed6AlgtJYhP29lxyphaaDIR8CGLv7bjAGHq
I0+TzcmIZAwi3vCDgWuUwP/V28QJ0X8tnksQ+vQo3zkc2izQrBDolWrBz6ZSwxAKEdktZnmIgxWX
JXjgnSfssDKV6GqYnyS0c5fdnW6sbp3EQJi+IIZLPieHscQ50r9ar/M95v/Ow7GzLx1iROAmnwED
xDmdz7zq9gN2Lu0upU2Qy4ctFVb8m+RIIktLuwO1z/3w2ThpTeYy7/cJeCsWNSk2QCL1/OapBad7
QmRwCwEPHvZYSqOqSw57CIFkFyaiPAgUPFj2hAuD9ER4ELIzf0gpdYcoz2KXkvaO4XNiConHPug0
mwhkzr54No5Yo9oJGCR1JLu/Uwp38I+1NqmWZBWRfIrn0uOZJew81gEsTEY1Oc9tqVniFqcWKwxE
/GZMzWIL2lX52Wk/ABWnZpQsZFfONTzsBO9rotSzffqXQ1CjiS6z2uNuCb4tcuI8hugTbEyMyQRi
+OyV4RnDCNhR2TsujMRsfQRA/NFcsCnS0FUjaazd9cXWq7WDFsIj2AcZqrWd0eWcq0Ioe4ALR8pE
SkoUGQXdj/sj6LQun91tDq91MfmG3SxX1u/jYbkhisgHCJszO2Zia4fQrP0CrLfTgPcXIJ607B68
QCs5sIWOc64nekEi7D9Lb8rvOgOcBt5ABkf3ZaIiVm5/7xlI38D/gO971aPjjamXiSg++bohE6Wv
/jHPfapc5nBGmVshp+8s7bwuxo/GtLF6Olpo3k5yi3O3eZeqN3iP9cQ4UjjoVUzio7iPyd/i68va
tl3XqkdQeL1zTsLH2aXDFnMNYmTxFN0oFo5Fp249ur8/iFcpuya8k3q65XLPujoair2k48ifVLqp
NNVYXxHSFpomR+qcAnmcwYyHb0b1CPNysojUJZPpmXlfQ5HxEQBpg13q4UuSH23WHeMi1AFQtYDU
JZiDGTn/yHtIPRzjaZ63SBpDorNG52NANFgo604zE1VqYZ1DXB5R1c/C09aWn9/4jgfDdljrO4DQ
AMHSCeLfV3f4uS6Xh98/z4sySSvCEH1O8lh1Y3HZBQduzh7v1gA6ub9Sq7XzrdErumd+2FMSB/dF
h7qj/7YVwqvc1Nyu2O9qLXs5yexKe1APNpWzRZK6rcF0mb71X9ujK50S7dcS2+1J8Q70Q7QVw7Dj
k1tgN73OvzN1z20juN9EssDnyzuSg+blqZJ0OwU98mRSGsWBbUhWxe84ArKH/CsC25CM588CFmjU
L4PFLhfUh1/+kr+3F5s7FhwngqaiPrM2YH6u2+v8VGuJ51hjkOYMmqUNP5bsetQuRHzWUVdNT2PN
/ZM3gUedfRKOknKHljJhv6DDXWtGyCl9/tRufi9Kn2RgFITCsfmFRwQJx8rzEYJkDD7urF7Tch49
hLgoAi4njwTn/oJkEDeeI1oD61q21nRrKYZ3dZOANBpD5/GJ3fCDNkxdM51WKqck3G3Xiuyfxge8
b2hYTxQThGtyJwNRmuLup8kY9NMnljWMHZ2rDY1n5ysbYYtijb2xNIn3pWO6XzhrKA9rc91P72jb
EMswGqf5w1nmjgP6/K4v5On2z3XvQgExCoYUfW1pbWCiCNV7zYDoyCEibkE3d9Y3DQsE5yqMNpPH
8UqeMkxbKZpmjYwFp49uFM6pogfL+U/AK7eiSZknOu6ndeIAuK1xUGuUMgJjTsPHXlrZ0aKPkQnT
OawoKU8DpRLISIqW9H3YRlHctifB1y7yDreY7gy18rMzy5Y+xjH11FNKoyKh0ywUerL5/m+Q2qkj
RX5g4S2ewEPz72LQMO0Xo8q/Csa1jXSIiPRSMLJU0SSKiE0g2NKVU5maVaIvnbTf6mPUedk9Avdu
mJ3s3EabZdtC67YNL4DlsYMRAApmAEhQDEFvpx8MhIDbsbVCwIFT/vSkxEl8CvZxytxR+i7Yijuk
GgzAKYpwXoJcL81DuhpSSJ6HJPjP0Kp1mz20NvEOQ3CkBc2OQS0KJjJup0naOF2ThQNVJwNuvZcO
tUxXId6p4lShBKO2FFlR0bplEFdhP0CYpQ9dZGKTG0rPl56jQKM6Cqi22AW8U4sp7ulYMeg8p1nH
pluEkpKAC+ng1DD0wRjV83Sp8cYlIRwoLRng1+17Qst3JwXYXDL0Y3pyazinYYsX87Zvy4jWn9K3
lkavulm/5m+Iazq40xZfb1Dux9dC6Z1pbQUZecYn3FVQy9J39EUYHg4q32g39usNqMZbEjuRTMi6
2PHhmW1XHd7kTovW9b7VbbKu/1QL32dGpKj7lJcqsSvMWpQuDc/OfkHqvMtVGFO3zSEC4jzGJ4b8
UERAsVZmMDnYt3DsXxhKxN1R7ZKaZ5mBk8AlvfWcJw9woblUp8ql0DZ9JANZgmZcr+LZ4TXUOzU/
dXOg5vDeQrHfLDxNf6bhEnpaEJkfifB85MN05nPEjbarNFYIiRCwtd9A5juiUdJrRhXLwCXydZR0
rKBtLzs1MZth1bofxWINWjUC4ku3iaJ2iMqWtutCv3ptHcXWjwbQMvLUiDabpVYo2Ak+IXtANvuJ
qqxUvwaRywqrGO9KwCXOqSXEtHQqPxIfZyR+1uxu7bCjuU6BV/AKw0YkRcEwhjA3kxxHByF+1r8Q
5qlF4TVz2sUeM4l6uUEqhhNKRomThtnFlmrmNB82zwso1XlPFWMl/Z0JvO0VZlBvM3ZeoRnDnqgd
V77oTiw5MfRTFMtNXaWpWmhuBR8wPLr1Kfi9if0oku/aNQFJKD2ANOHheQMIDVfExQ2LD5SDEWkZ
RiZI3fa8d2QzAUogBb1ODj08A0ESr6WhNFFnXdIt6f3xnjqM+Rp934/TpGkNNS6+kv/ab3cTdSSj
sbKoP8ig5USswk2Bcu4Bh5+RdslXZ1a3eBkrIF6ut4BbBKt/3bNwFJVX8MksalhKxJSdk3w7tGgB
bp6tw09lOseLYeE4A/QRoC2Mt3ou+PnTgziczGYRQTynJOGOmQMcbdk5Q8Z1xuxk6uBEyFQkFu1+
PqmZJk0PEApUJRk6nhaiWJKhJilau6CpgBJbo90B9U26rtsvhUdxSjTskIZeODfTKs3gcxVmZ7O9
PxE1BcNlUzUE9A447eL0RWwkN4pCV+tFZXlIFvWWhlTipUHyk5Eh5uZOOVud3m1x8CfH5LglTLEY
s1Oa2wnEGb/zRIfbWSPiooAx7DA3soVYQi6rEg/iANm0ykVAYt/0h5YLIvH49dq82pEgI59PDctb
WeokFcmji/nQB5wXvCeGZXOwUHLR6iyHQX7R1Qsuj9YXbCrLOpZYczQxCPOlggzzylkbukhMDOyE
t+bVA/O+Tutx2WtE1xI1oJd42uUc+M40P8KctG/DmoH8k6WmErDMIapUDG/cRTHM1EuUgCiEmvht
JDbywO/Im8AqCSu40OjRhV7Z2QSmbe43E/wfMXxO6IzRsWyYxkKz28ol+/WcEjaDOvQtmrAZBuiB
cJdPnpbfrdS84dQIFtQPOGNiGK2Wq2jCS0ob79etJykJ9WISWKmAluWPO6tFeoJhNeTMEs3JD/S4
ytNk3FZ684bbG7VCllIOaV6QdZTqIdCsu6RetCuepnW17OtkPkhXz344ZlbnRz1OESY5zMYposYa
d537Lw9bhWlBaXqTFhPikGFq/AG4jerAJv5h4p4aT6c53vYGiK/hvAztQ6A8f48iJ8J1sbTbWzo2
bef5sfizDRgg4YSs21LP2QKhxHWV20L574V9DHtdkcHGHcoHTV7HBj1pRczQzbu6gS7EgB8SCnPc
IyCXR/tMqQtQRG0svyYXsLaPjYzliX6668rWNN/rw4tsQqAPSvaU4vbXNQTgycMwzSKxAS/gkLc8
wlfZkCSNeGi+8ilRZX0g7BQKF9x318mMQF38ka4XbmEHwyY+GgoAv3YtBUqQZiZaVM3K1lwRwVJt
yrwoRrQEW3MkuWHgUHrWVIA2gLSoOMeQW8KgNmrtzyMfEGUj3BgfLv6nIVS9RxyQ1dl2KWBDoknz
d06iSeg/0npbRYLnee3mKOoAF4csoZFY/WXZfhaiS7MbFrmOVB+GWvK9A0ihesFibtzGPNmoY4Yh
TtqiPn4Lhm+Igtapayt27qZxjVRIws7f2xiehP5VVaC6o8jnzkkQ45aLNEGBRmRbuzPlPAoENrn/
sxtHim2QWLCtcT9TCHQAVoIQJDCzFS15hJZ3p9aMua6LiVJ+NFa7PKoU3ttMbIKuUL+bDXG0OR1P
KZGE9exA/aqgHgnr5tuIESp3oRaIkSLEnySCxEUgZ9DwP+iMgw1pqvFRAlEgvf5V8xiRfhZmpvmM
P2y1x2FYJUszBVU75tq3PD3+BVOo88zg37MaP7XOUsChQDQ1o3rLYor0AKXkNdhr5+x7Zg0m/uGq
OFzEf7V0PiSushng+yQStTXXc/F5NxRExIMMNkVlFVVe0OM9VFb3OQyAO6LOaiN70cd+1T4rLzv+
IGLbmvqOHs8A5Nb5kU+VGjDl+yPVs16PyFHNXdsghq4zLhrLUX8llztuEPnKs3Nw9f4hNMa/QUb3
GqskW07SGgxMHJS6nU6db496hnZ0RJHSapIs+k9yj9urqEV1S/266Z2b4AsX5LNacgKP0LUcLHY9
nO5zbzsV6ZTFVDCVa8xTxn9XVBGlvQGdXadCylzbnOlx4nsZOHo5bsnhC91RgBST7nlzfhtpMj33
VRePX0P99WwsqEKR2ukTQNyhxQob4M8HEGUkV7mAbMBdBS6vrEzUyi5uR6novBERfyiX9nodDo+F
yn9wDuAgx54Tl51XhRvGfAPnCJ22dAVQy6dsLQrVnlGHG1yuGuA5ju8cjnGtS4nM/PrLtsOGOWMn
Plv7qJj34UHXRMFVOOAIvCG96+2seVPLufbThiIiGpRp4hNTrbL6hESgnP0A4ocFEyhOlSBH6mX6
LS+dsHMn1RvQOd6rGVqiU8pA6PJDlIls/RMnGkXVbOcn7PuD7qe5QLTG2jibnpmo2zyJvjEza96g
7R39qKwJE4YTit/8bIO1aNTAjb3BpKGfrSR+L9M3R9MGoC/ARKz7pkhjdJ/nBz5udFPMRzR2/YZ+
pmK5UYymwnhJadrLINKem1jdANRcolXQ8H1ex6PTdi4kX0/rSSaWQxU6PBfXKgmnJ1WPjBtK7JZh
FRB8hxxJDU35NQReWf2/Px7EDF/1FYJE9iwWMVEiigM2OjlAr/ayFDaY2kxYhw2c2Cgj7VaR0qWG
5vUN6iLgpfd5CSELM6FSb72O1vC8uTIlV5TqxyYObpm1oHDIoJhSxPPNbk3ZH+xHWTNKI3VlnOVj
S/wc2TIsweoBtQyHTMEK6jQbNIQ7vEOo75zqj1l44GdLTIDo00TDTr6F99ak37CPbGkrLIqr04P3
S2JvjoU+lcdwNiNYBg7U6wWySrH7uBC+Fy93DH4JHQ21Ok/VGEYW+MYQHxhcL1rIoBzibT+UahxN
6fYTYkeMlkmd15SC1rg8rRq/fRf5COFRUYyTEhrEAcr5WGs2j58P/xQKHc9nw5Ox6qoix/CWzBmZ
14Pfti7Yp2zTPcJg2eXGNdazsvvm194o+QHLFAkYjBqGA+Bs8ja8+C5mWCwyd0z5oLbvNuH7GWPv
272I4nuP6OihhLeG+8TnNMgQX9eYqVZynf4GAl6G4SDV3BLQToj5YeT1pX5is4glopqjzcY40WDI
QElq7s1iBkHyH0ee3Kmqy3MooNNBU0jk+Cm9BFZYmBkGLUftQwZMzOeO99mn3L3petM5nGYZyILS
bMCuYQCaoC4RfQeOuyxaLcSIHc9Yt3xewY8g634kwTG71vokSwkxO3Efc2H9f1soO0UZjM1BjBSX
YIASxiraL3NSr5Et0MCpkTJ8WLGQXKD2TNvxa2YR6tQKq8+TJcyXfGuxrVIWi+85gVGPncHsBy2h
Adp4Z3cWBMPfjI5e8PSjOW8HyEq8x9zI/ta4qxucgtUPfh/aqpCpbYZeiUpk2AzuJXlq4VDDDrTa
ry1QkR8qo46zz35WdfTAgDU0f92wqjntmbc2pvvk/iY7jfkXdolfn3v9KlQfm2PA2FXL/d3cVnQp
9VwC7MegTvMBIprZzN5+FSCWmMFLI+MuMOweB5uk/Z313AtwhJdZkuvgJGQqd7EI6gj3hI+RAi1P
YfUPbr9qwJ28b7QRNat/S+Ky4z8vkXkx9dHf+xw5PwKB2gNNIE/fSU9kEecQu7ZulEF7ChJmlubu
3GPc8GfeKzfOtc1b3Bq+kqA5v+cJ+4gTTpfmv/ng1VEfovbv9GiNQZqXJWF8zSZiOwKjD/ayhoGf
n2G1ff13WbrGjvoU/QSbU2kpqACanM/HZWmobaL4HQiL0UoI2uMtFKRVOHq2DJYyC4GKv+ooTeyH
9/3eMHG3ODJp/1XMFdyC6JfPIflW1atx8+XQH3RJzK4UaJpMPsL/K20J25MMOAvgSyEAe1hhdxzk
n9HN8Z7yjJI80G2K9aBV8ZKliriaa7Kezv71dTm2qr7c6IAQybIX+AIaNaNLSbT+2EpEHTuBYLO7
sI2903A6IibMcnJ0+42oqRF1tzobnWbDxK+NeoMYnaJt+SzylMZdd47wTMOH8DvYqnrZLKiezdDG
pojFJqwka0ZFpgXAEFZ6ZzwkKz8iCm5MC47G84nQP+YNvjQb7zZz57ZiIzvw1y019lZszfdP3seP
YM95UGnEbSg6395Kil20j7Tp552jksKTSZ+VS1aSHCije/2FAhiNtcUN0C8CkCQXzDEazFknEEja
LaT0ye1fVkqcLLbVzvhf/Wk1AMxf4YjrRGddGWCNxMrEfQqjC3PZtyqIQnoWFVjCPCUvggn0uyMH
bwaSS7XpTx+Rwtvg8SDKDVsbnIUDFkhJNb3QcOxGomLx+dTTNPlVaR/ZooTucp2ZTGKJrxOPEV02
tPxx9zbOomamEaayjd2xEoyt0DLxeDBmrHiOFO38QGFFSHhS4Y5swNL7NqFG4cyrHgywBSFV5c5M
MG1jDK8pOCDkokq7K/cSG36CV+ff9SOqD9MZBWEC+6KjngkfKThf/V2ZN8qiLT3+C9LGKpeTu4V+
OCkRrxvHoQX8NS1dt2P/Hedq9ueHjrvUJaks6f1b0hWogKRTAbdcC1Z9lhK9fYSqFiFzemO6+Oms
B2H+CuETOXHlJZpeNj0jKH2j7bpTvDqSeJziw9crpzNFSRQbNtN+5HHVwUKp9eO4+dgI1AkuSI5E
JGHkpHiTv8Oua2/di6EoNYtYltRtojcJFx6QnvfddvEGu/fbpIOnHWNURxoR3z0p22IbFdMS8YoH
lQJOXRiKWL1mJuP2Kj+3dTALO0Q/9j2Cm7mczgHya3u/Z+caXvWwYzWq3mShi9HMVm7SXaZiCfB2
kFqEAJafVAE+Zp/NjNoRjYPt/sfWjOQ08sdHJ+rq/880IBxDYYqoeWPJivaFJHAH42llHNluWNaq
g7uaEIDhJce+SqnAaa7apjbDu6MMjUfsA0ONa9RcM/LDLZoFvVDRUHdY65ZlxGcf5zthUMqvs4nm
AOwEND3+/UllpTgP2Jqiu4HCu7Sj28PKfuvrfCtKq6ZX37QfOFzyDeDLiazY0f7SxRMa0SVNmHIn
MvCgUoCZr32QJEgMjHtAsySu/qbuoooxNRUYa3AJ2qMs75+ZkkkYKG04Uhol4NcXZP9JPbUnMgFH
Tx/XouSq3gYk4YoM1AUpwwlLXXBFAeP0dR4iZZI2DOJdV15H/FShyn/wR7hj9T4MeZGQvG++U3LX
3FKBCIrWLtX40MgAg5u0P1Tc7uTL0hO0s+30kNoOEO2W34K6yJFoXahl+PC/Kwob+2cBdHZipt72
kMVzunMK2CpTFJMDiAkaIAfctNrrzqytkVucjgyWyosCEzK6Xh2Nq+HqIkXCprYrZ/TcX6pTO3zW
mP3VWRQoAutG8ox9+6wuH3Qmy061H5eMjXNioD23txqScbJD8YhRtjilHF6pndtYK/6td2Jp0Q9F
Yn4oaG+6Lk0pebleWFUdoY1kqPQdFB3l8YoTpOSdSX63T5Mpkimy0P0rFMZePgYJHmrAdyvGvACX
d0W8U4SUbsCOASUOS1UfXTsp4NoM32Za5VCfK1hynGb7WPcsBzhyW2bd+FO8TiuCTLmtD9dcW2dW
h6yBfqdetteQwN1mvKEPDprT3T5F7SMKxGOz0YxsKUTG9HfK1GtL5t5ri1VtHt67T9+OSMgLQt4Y
7hCrFwOaAGgsYVt2V6b8p5BqeBcUzXVaxFXPI323l7KpleUIveq/7MbPVzoQwXTEAmogGg4vifrG
Hp2qRjnNwohth53tr09fUeghtZOmg+sRGt8lGJwbt8x9iDF+Ve5wqsedIk8FhZ20xPGDHjEZoh4w
Vfu5dG4BBs1tiPw0OU9H0BQNG6ZmcReBWO85mdAa8vJRynUexgEt+3hi2XEqlCi6SCDck1t7fo9D
qIDaLrNZ2zyHokiG1gn63MmVXKKKMgW93ohOzXUASRzlb2reYuAwhhe3OVIk1nxP/bNFTg3UcneB
MGIrLPg8oJBVwBnebshM2MwBrxFlEBojnZRuxlgZ47J8QAblMRI3fkEi9Zy1in7OEZoWCAg379EU
PkXfu7+LiTBKYREy73oLdDAq9laragdW7auk3hPto7EyYgkTvmR1ZaJrZhOx36X2ODg9upOtt2Cg
FmUx9GdxgqIkYVPGHeqIK8UVMh9G+m4vRL6H7nsbkK9w/G0xmfwGrjG8EYgfvSPrIaPM0fgbeRR7
7w/ZQ9ESWttThZfGv5pOjk+KPucbsezBGcwrDb5z4Oc/j82FJSE0Oaf5eyEJI6dxH28db18/8jo1
5QogwynsM7x2KD9dldcvEfYLhPezK8ADmQJLczGWlj9yWNJbNhMpqbmeJKWBGWVk+dTSFHxaDsbo
KCE+C2CnXK52kI61t0h0wX38p3zSFJRk8a1o4+mvmwYeHymKuti4/Vb+nf6e19jXdheAv4Ib6M6w
9X/maiRWybCeczwuA4m7zq0z4+aOsouf0G1oi5QgY1ovBXdycYeHN4BZBooJ5hDmlJCokfFTk7cT
pJqLaHozJ6H9A2LeN02G4p8x5Y2YoeZCAr6hyZidGRhU7lNkFTgU+FCuL4d3dvzCwyX85P8kwAjj
rDz/RLvcWfbgFBvOjswsB8b2JQLYmEv4lx6Qw9b/xxRKCiDieQxhUEtjkCCbsOAI/UiBA5Tn+fAw
XBOn2+7+e3pIzNa0uW+ZGdH0DV//9ZM/5ChrTgk6okbYo2jclvPW1GBKXALJlVhiaVg0LuK5c5RO
AIaJd3eqsb2z98z7ZNtmckF6t04SHvwJNHyTT9xh7cQ2ZSgwqKNzatU0mHe5S8qhWowOFKulyeMC
2UZX7Ih35YjmEFYHH4OrYBetqPNpZQ/6sA/kPmcHFaPWdSRt6M4XXE95TnSJ+yl6lQWkVCWlhf3o
hr4hKSWgDejmYvqhNwh6dTqZ7/CjhQysQ/70WQojjAcNeqTBcr0Iu3z1zzUQk7etpgoWxiHYJsng
RFGm9MfaSuCPRRE/ZiByp1QAGpsp2Km6zIt25NYXlkj2xXfHnDf09WEFiFUkC1h/l/uG+1rKyjvz
7BFJIiNETz8Vb6H3xocjSuDteKk7xoQqQel0bQaRYNhqe4DrDa6BIWO9ZXOJmjB9lLB62MSjj1y+
HsBh5e7AgXKS3Oqt3GFp4+MXPYdVmrlXQ6vhFFkVFmmCIIZ3KUUppn8vIOyjfluXCfJ+nB4jda7i
tlrDgX3qGBdhjVoN+sHUzN/bfT0CPvO1vVyPMnGxzsIeAmCAZy2tWWAxyBjLYbNMGh7iCahJ1AAA
3ZMYoJqnAYfHjMW0eXAd3goR4wQ6tZRka9tJObfo5zafB7MJ+VsdvEJzj4Hnb8+GHj1BXCsDbfyH
QichVP3LliZ3nLn+cKkh7p9ivMqqgNcp6NM+TMwZI3kKfLtP7g8cbWm95ddszlpCHXYEwyrrr1eD
F7+fFRjm0wLqaKhRB92pZzWDemGwxoYz+UUomXwgkLmkgEMhORXI9R4MquDsLig+njEKokCetKeh
0TBqtXMZuC7mH6/+/4zAcvPm7XXoXyaGHscJMvyCP8E/zIIY+3BN2tdOVDaOJtcvKqX214/VKSR2
w8zEsF7OPseg9slQV+K3X5W8eYR2SuYkQ6bwrr0uHhB4fkbRpQThfLvqmmo5eWbYFcJXJ3GnKvlw
cl/n9WkxkyGXOZQ8ZEmoFPLl2wxbhV/5eq0ZhxKboz+LmGP1llMu1poLCE9pRMmKOFA52bguAdwz
YExxCEwsi04AFQWl2fcLHRIv3dO5lZclsXapHSHCFaJgrVqGMqH3LDl6himjFL5GjPEoOGzFWWvr
RJUugoI6SNArJnpNl8SCb44RSTsHhxsK/xNIYH4NjdhpO1s3GCDHCoeHoJ/RBltdJtkeqB5xjh9s
zFTpKpvm9LQa7ima9PY+PokayYcOeBKEfr09FUSl/CPM09tpUA0w4NwZsHPaXqWGMIcQzFXh78vZ
S0vcvfh3enUpDR9DVjCEiHIikDfsafPbA0sVd0M1AeqzBsdrXYLBz/lyz96KdA4LF7k41j183+0V
zmuSnlSv5n6BsS2CBMMkaHyHbrBtE0fFuoj7CXkIxw0rcVN+YdHr/zYSkh9fR1/OY705VxmX3Vil
vD3zKuEJTtwTUSImLzR+3UyeT79WlVceRn5Tk3gc56V7B7t9JWW/MeVqu+WO/CPFvucRdXShykDm
FaFNgTHIScDX6d+0ne+WULww2yfsHu+ECPvEOFNsMcfGMYd1ZxHG0tZSQq0bzkx+uyHTedJiP/Q+
MOTptz3yiLGX7ZOw1WuCWjpJnUajjXmW0RpqbPZESdfiVvimvuykvBdixorW+JWqPsGMn0uxwx3b
bJpYILHCNtKzqAsZc5nk++Ea22ipULeUgufodx9ZN2SS8cJMUCql3ZQVouTTjrVsFirrPYReoKm/
y6Ow8swrVIlHXBgB8ns4TUSbfjduk/Z+HPkX5FwxahxDHZYJ+QMlp1RsQnlk2HpQkR0VV+mjS7QS
wdcN6yn56YGX+tNuILFrYDk1863tK23JekSG56wZBvkuAad9Lp2VEDIhsHq167LiWLrVuvbKQ16B
Dpx8wCw45h4fmxtc3sIiSPmGWUptYlLuYEEf+dtnO64vQa2wJ8BEdjIICKmsvmLRUVeG6Q3XS/ix
NNL1JuteELn7j5rKXdaAvZvDcG9piZbVl/gwuD6/wWQX+NMrVwqoIzpv9oePIZvdCOyyvnnYnn/m
fT6ti64Hcr8RV+lyrzbGZQzPpc0M1oj1pNY6SZNDvT6R30Bv+sBxkVVS9WQvlR9/O6vS97oecZij
+QpEVAK9eA25SB8s2bIyqJk8in8DHBfb8XRYn1SMacungR6hZ+Zk1gtqufIA0G/XJg3YUc8qMium
pv2EMaUQkGbsPn5nhrFPiP/4/3BxB3jz365TUzm8p5sBvYTg4QNyYqvQza5Ev6pUz2ZPOKTTCfmk
byP4T37DZ9XF/gDi0RHVWYILzkw1XuGi2YIStMBc8a7lHO9Yyv6r2t7G0uCklcda49YyYVoMXW7K
hXHump03YD96k0cjfnd+ZaPM9WECHTSxhS1cdtEOC9nNRtvhqYaegEECOsq/ZC6ChgBwWAzq14RC
qTczhIixqUVp559shetA5G5ioWhvVwAdf3JHdHUeZ/JSD9GAcS1sQ0abyyfeiFiu+KcuD11t93Ds
bFPMZzc54lnNtbdAxiBIdCZ14TaPggvcn0SO71njUJiQRiiQkUdh93POWOy9Gy4C5lTCviNrOv77
BiePrcsA7Ot6+e8BSzQkfa1dn5cGwOJwIro5wmvb2jreMEL4tjLryFFGg3dwnHDcPVCCOxLG6D71
UrBSWz6nyNGfGBcrJ8stuMKS6TYGRua0c3WpgvbJ3tx4GsuaD7YKO+4Ls9ePzd3/VjW3PVm3aXqd
+2Q+DCMdfqTKQOgO8+xJWsSgm/VnzK/110KFNVCYV0dtr5qjHEHeQwYAhZrbMOfbMcvu8trGIKAJ
s3IGHlLK/133aSkgbrWTWpyJQ/J35W0xaIuKpo2KvMzBStx+wk1hYAwTm59gDVHfP5jyG2dmBmZ9
Vsk0kLsIl4Mm3I6Erk7ohBFGMYG3bLGXw6cYQ+nzHl0Ocpor8De1dwZ3X8mDaozrBKad7C9dnDZj
SGxQDZMU2yWvNGiUpxzFMYQVz4ONWZ9pb0CGC/5acg5lZIE4kmR7MxtivPS7s5VSIqe8qmw2CaKx
avmXKrVxbRzzQK7Gblete0RDmbs84ittEbqVdp0XCuR+HQ72s3Ru2I6W8gCYB2Wgymmxl1BIs+a5
0i78hvsSAM8Ku6lGr7piBT9jqbahDa6ER/ClnaRm7kbabYbI4ZiraPYHaAmkcAmWMMwcABP59Q9l
bmQIRqcjoBKnCZhJAEh5GocwpOxLT2+Vc5+GqJ0TyqFj+fbb4rDQfYEsDssDw5Af7xwIqkEcTW0y
O8+o2FyTHOoddusnlZI/BFD8p9JRMDis63VyizTQKu4KvnZcc08kB1Zow9TzW9hJITYw/y2Q9umS
o2I/dppMrpp756WIJDEv91/v9pfb/HFqL4V/Lfzsfr/wbhlInXMSuja22AW6OHk0snJAgzmknQUm
lcwQQP44va77Nvs9+nvfVBmr95wLOQziveX5c1HlkwvzG7JFE415gEAVCyJoc6aaCI3KicREvmpa
qQNyShaa1be5lFjaOMz0o8syvwtlLkiBbCK6PifK3z/DHY/v5gVjH7Ja3EA3hF4y/Vg16imtKdZt
KZ46GtNbfTD03AsGfe4Hh0NvaZsf+/lUMMUGCZygQv0XYDQ8ZpDSuSxs6nIrtNHgwWSJEBFuLyIB
rguvsprhy/11E+uGcUK7f8wgNrk9/btuma9oPi/M7Fwx+HwuMJulR+OLw+a3bYhRTD32mmipDEE1
5EErIYD6mjZ/t0iIng7CaCpRGLq0J5mZld1p3wxo8Hloh1VuH01usIlrBdbfngaQKQHTOt4J7bNb
4Cbhof1nuO1+2+awiKF19Zek1SQcdTAxbtejfl7U4DuqN4T6BTtrtRlLR5PhCJKBFQi+wA/5O6ub
jWaPDIdSDQt7lAwNYG5wN+yNWquSeRpElsieKWklRvCEyHy9E6ysEy6C1UlIlhnqFf/zRS9PilLG
uOOhVXJsdP23c8Da97p0ZM6WXt/9H1JE4IXLFfjOSbc8vpm66bWDTN/3++u9hKFxOGrQ/jzO3Z21
jwYAZtXX6BQGvdFtr2DAu+Q8PM11PdtXb/wPj3178y3KASvBggOffLGelpKUKvhrXWt6dOjBBrQX
/5+rhsQ6K0IXtqNLZvzUYY407c2HaNaYK7V7FJ2cOTIiFV12w1rBxBDhDMnP2f8KBtdcWbzwsfGC
U9PbkANJ4VPPV6Eki5vCFC95RD4y9gPw+9pTkwUxSCid9HiEoS1n+bUHctlgPk6qLbCTUmr+DNrJ
BZ6UER1TFKVhlZ3HcE1nZqdWVKteE2DUvBV4WLZi5by4EtDLr4Ol60mKLOYlKJSUrLzma+Y3NXv/
sTy3V+oWx7Sh7R+n/ukZtznlYjJZ4NfWuPU8Bpvc4WDeiFB/KL+U7jG6B9avOR/+eiJnu9G2AWs5
5p0LrGNTvFVKsQKG2ub04nW9gTu/fbmkuAfQ5J4QGnTqaDXXAhdrImfHRYVSl7WO/+J3OnFGZU+F
QFpEwly1MwowafpHZoVjlpWX6RZhfTFtSYoi0cSqDN/ZxJDOXsXjAnFDPt4aiTW6MwNDSjL8NPuV
Gzj+p32+wa+0iuY2beTaNUMns1IQ/3Xy2RG5BJgDSb5EdN5vU/wGLztwtQal5fyC0wSJzZmR6f0L
YnhbiTRerJkb292mGSVJ1rkreHGOfFgWnAaAoYd3mVj+LdPS/cg6l75XkSs2Sm3MvvgO3d0W1Xy8
Pm9Hf8ge6wivnZWxjrd3X4i45KrcasFjaquPLmq9LCFmAzCyWcBXkQCeLdDvDibznqgArLQfQX+A
EoF763AgKPFRPhwPakjQbBoSW4lO8dAkeoLPgRVgUzf2FzFLbs38XW/mCdFhIZH3SC1ngz5h8JPn
cGSHsZ0+O5qxYTXqh1BcNWzVlTlvkB1eVf8nkgFRP4JdGuOUuPi6eUeLP+4Mpz9SA9mZKDmpNL42
NjDWrpB5KKCVQhKA3KpRH/Qflq1Y5/VmmkU3BFEw+k+1u5NBAL0ZCyhnBvyqdxMV3qD+p0YTzM5k
TDKoMSWX5S6gqL5eR/PIaRWVSpgSl1tw9J4o5+lBjEubYH8ZPt5tu6ZGqFJy1oRzb7+nj4GJcYr4
pe4k5OIZY5396COkSw8m//3yKv7Yg5lbpSQM0+wJSH3oT6HKFCfZEcq1TkN9RyWgObUmSbBgtoJ0
VuULP09hBBQKoLhMncWk+b7DKTHO2gtaVVWIsUgGYqsPGDAx+lLsUSVyzOVZ43Tp/+eLOF9H+qmD
l9uhDNwQxxkwohC5ARPtlJD3CPdzcYby8LrCP70xkeTz4O5ytEBL4gHfDF81cUp7z2m7axK+EPNq
/a2Tiqi8goFbmM26LIrZ7TPQg4dR5ae6CevLGO/8VX62iAW5xHEiPOaItjl85mHPeuG3/gVehNHK
1P31BqULU/mV+LsT5SUWfitBBW0qxytmj6YHnjgsrKIsm2jD6lzk9v6OKcZSach1WOwhpADSu4Iq
CFpg5cFg9NoOh0sQfd+1vJ9PRR14RmP+/+4aRk9DnV941ZsVcF4mD8sMaUVaLqv48aWsd0zIQw7Y
ddYB2lgLe50WgSSMDwDwanrEXm1OfXJdx6HVB9PwHzYvd8f3FRHZtTUj3vxkF+ZE445VLZfLQ8Oj
/ILcrZXBUotYAvKqTFAG4YzfLboh9VNdsGaMqA0QkZq/+VkOvgoki3As97oMAgoBY0sWc850OvjU
urADTDPdevC6LaQAwzuJGqzOtO2qbbHDjRzV8Sr41ef1Ri0brw/yUsJ478Xl6Ek1ZFicr0eTaFu7
pxld31msuJLWFh6yjtyi03Pk8H9zf/XZ1t+98fIxPZRq70vuEOxtkknjNjAZKPgcCZxrHCdZsrQz
KBI0VZwNq7fHkoJnvV8KhW2rpkDulgQVJZDzcmgwMJfpZ7LaFkSxtsj1dxo5uQlrFhcOIIuYxbzq
TU3Heug6Nfxu85a9S3QXNYSXgURJDIX1bcwC23PZsI4m/oSetNs3r87nvDDE2U8wlBGiD9Oh2GOM
UVJJ8eqjqqZ14di4xnaP7xbgsnJdyKeqjczhD424eFRCscLFyW6lP+TKjuXGROqq+otGCAsVKAAM
Ar/7/vslB12h785rY7N1M6ScalIcJgk/g9KfF1l+OhbObIp35w9GRv5nZWX354vdOWxvXjroez/e
CmXfAxK0njNkjXAA0s6uskwcicfjEhyyLOB77dI5ZzIk7Y4T1lHUcv9e2neh762b8WkDGnCJHqQl
wWDH3N103y6qP3q+4FG7z1o4oFT3nO8dG6lZ4VevziGjuOBVyy2JgezANjERlZxCfl9t+rihATos
kBaBVBBn8idAycHKdwGQzevyjcYQQkd3Xt/3qQulc5f+5/tK7QrQQEmu5zzbSCndtOEyoXosDQRm
MmLoazNSZDBsBt6YDEm8vE4R0NA3UeC8X1s7HK8bTC/hQuA7a4JG4pyefZwXAn8VnZw9JhsMQJNR
pFDhvljtY9nlmsx1zVOtv0glKScLgwNDdPmqNO9wn6fuI98bDfliHavG8slPyq9I+h/VBMunYZ4X
/F4dO6jT+SLtwpv4nbU0qtTCHYHU7HnqSlD08DmnDbpg7NYQDaHNeCmf8SVeiL9hv4N+YbVZMtCV
yfiN6Cf7KB1DAn5bczggcu67TvuPo0RJr9crFsQ8Y5Z8u/6w+exGzWFjauWL0skzi8fzpRJTvEtD
fV1NlGYgdn2FsrzNwY3HEU6r3NXZgfuimEqYGTERo762SjpWPrnCQWyVnDzMuZOoWvnJ3f0+ixJ6
UeQH/SFkvWxYrBol3otI3F+YxnPEOe3eQ1XWYM6rgQmqh2yRhpPPno/4jPyrSL7htDsrlecNqcz9
UJP3o9K5Lg21FhPREzzJQIsSoNgwln0K50FaX8Bc8RUyPNdpW2fiUsyIuGu7UKG6oazpHfxPo8YM
17rDUm3XP5c9JhOSCcu4DKTW99NmwynN7rGxYfZ+CWzXkkWY1JTWqME6dEZ1oxgYySGZuDudambw
Q4Raj9Z/TLVPA9CpHKlYSDJi4Y82MHC537pQIgV1fbUN0IQCZTJcv9gcMJTeQGkeJCy00QB8SP5t
whyPLMKMj2gYqQgLFRp+910H5u3NxjS/HtGIvXRvqfTr7mh/gCpbb47c23YiU2wmwS17+1dmw0yg
gJ7kH6bB6O94sRjDDeTlWMLVbJHzQ5CcbmZmsuuvgZ0hJzkmAiRrNva6IJE3t+4WJdyld8fDvvg2
va+NuNoakuRKvU4yj6HmRaMgM6M79bPtMqVfNng1YARWNW7ekrQtyxYuZngDbtYxI2tQVJpMjIs1
sW6xoGpf62tgp2etcaaRjP4dL734wb5+klmSEzsYIDjY++jRquy7lX3nuoOMB/+lByeLneCZQC5A
mWXgCQkP219ifkeDiWkM4hl+uMwijehTQZyJa8VffWV3powxRM/a5L7hvl7bm/9nkiifJVKdTMCP
VvS3xdRxhgKo/z5h3IAYNQIXomjBqFluS1Po+fvqfXJJU7R8yZHJLFqk5+CW9As8840hnEYj6UcR
t5/NmBJjolPgawi5gilvYwhfGKjURKoed0A1dm+qX6lLXSwnvlBab6i3X76kS/QQJ17KtX7X2Xjx
kLDg81OTkTAEAhyzCyqqjHbwE2cjbA95XxQwAxMkt9GLruARJZ+Ln7mWVyoR63UNVTu1NmLWySVT
tmanQUFT4X08/jwsfzGVLHcx7LxYG1mtnHQztBPVvJ3KUFrfFngAT1VAn5lpHrk1p4h12Jfk7+QV
jFBIF0ITwROy4nAryguZH5RzsaHLTzg4OiIqJgKF8OU+Yqz79CLMMC5EZ86hmoBJnxAyS8VPnCvp
Rv1wpAfEcX+rUNxsAR44eHs390iq6a6lkuqY9D8qbIZUDDuOJ1vCEg0hmryamIa20TuRW7N7xam7
VEkUXBjTzHTIBQP7FOl26IgAWvhyIxvL2a8WUUtLETsrBw/e8vontl8prvOl854t2JVXKLm7sdYb
mBWngDP8qIm0XtGbLlDvLXxgqf+odljVGnWMB+8T03+xe8NP/sWFuFnwjhmRc5VLhPKFIBqCtBL0
DJ6i8Y1DmeIK/c7wnGJPAoen5o9FSOFdRKHJjfymg3cJRM+2R4vTjAZqQ/ax5MZJc/v+iZbzJzes
bOZ0AqyEdkX9mnj5lMx+mIWvfwtkOPP0CELGUw7ZZoCt9aXWSR59rpMWeZPm1mzAyxwP08KjfiXz
o/cuEgZlDyf5U5SELrJk3ihmZIk2AcvZEqK9BdhKrtegpwp4PTkU4tqYogIW6p8UNcoALh6nIKMW
RVIOp4UouLDpn5nxENuCYiqwbpwYUBN+mzNMV8q3wJYUnfMGBOK5plw1FqK2ylvncSljoOikfnmD
FvXYED7hm9QrLaSvTuCX0ORN5dFmX4Tp/aPx1uzhKeesqxuagulMM5FAVS2X/0e0RbCPJkN/OPTI
hKGtLWs6A40+yhCnJdWeJnPJ6o+in8pX7MWMdrj9ZSKVIIaUsx59kh8pUMsg9FEmwX7vUOWKilna
RL1aKoJohpG+kuXKAIEMscek1N+49DHDeKawqVg+LWnjD4DEAPGZqRqmh8dXH2KnCbFke2qfP01z
4ck13CRhoa/ZIQoiBBIBpUAPD6n6lssPhEdhp7kpyr+y99Dst1xLaOfZmDBG+YeVntKgfZu4ayC+
wP9d3+AfpH/VVcaIgYZRMyQPjXCVQ0janVs4isCs8L2GBAbISZMeqwu5OcdTBP42c1r4YJnaCe6H
CRx8r2Y+6kA8rPzyNJkP+s3wSGKtzQNAA9ZkdCY4s4ombtnJFczvh2Fnpwr39RcRNYg9HHnfkZsT
LhDTi3gcICK0uDO58rG7wW27HbfP6ghUguFHmHnHiJHlHCqb2yxIWK522T1qq1Ps2Ji/tcXG8VNf
1m0N3JZlc+UEGZU1wynZKYRrHEUMCxiEFMGVBQtZDfrxcCVaX66yRNc+cR1C6kowOgbT4Mk0Bfok
1H6DwfDHapcqdAqGz3HzVQdBbVq5vfewC/YRLedcjbHEKxGfrgOynRAxds9p1XScQg1J69MJwePV
DMFoZuaXv6VDbjImPg4JzJAyuaNJnwiHbeL6m6hOm23fy+wYGdAzkpffGV5fM+5SZcyJNWvDwFaq
rF9mg6Dw7IkGWq95T8wocbz/CRiWqqEFlt4+dDgvUjN6H5Ir0GREw/6rIvD3AxANeuA+mbfq+7AN
nZM5nSluxpXVHH1oWRAwlRU4p++5Bx0XYJDau8CnLwUlXIZL8HJBSZH3c7tI43EE9KNK1Qvzw8yD
PQYgJdIVIlMOuKEeIsHpIlg7VZITYeDv/XmVyIkwP3xuPxg1a3wsWmsqZM55YOr9WByGgYYCerHJ
4TMckV7LQokUk7OLPiSkLczdUy/ij5oXAhNfohVnsxRQhbUsGb1gDdN5MZklsCP4X4p3qCem3VaJ
Q8ppmu9AwrmBufhW0RRkESkVOWdh6iUCH6f6Fx9kUdOJJIxGSoBhXHZJ1a64gVz9o0PMpYyB77SQ
zEvZS2onRlyQXLDBpVF6joPSovVxLwl52pua7MrxtSzL1OSrgECQN5S59qE3uby7Kmsr8BpicbuB
HP97ku1i0Dq0z1GZGkCzvlXYOX8JqpPDtCPRfnMXp1GhmVOf83Vmkxl9gFFaaM6ur2XG1ozi+RmE
plDQVLBdHYSzWVtWFX778t2Ue6WfZHLIh8egfW9DyMipUMl1elxxm3MwZHOLQWmxGEtrUHKZSZHS
vc2LgUppO/Xy+PEwNdFFodDOOQD+JCHuQ4ROqzhA7NWa4n6gqXCJsb0nHDecEyovmqQUtPv+wCe/
IJ4AG5FNZ/VOurx3iL26G09uJrYImk4z+Xlj9iq/D0BYhUkHGyqPBEqUOIiBR2krAJVuUE6Dm+aG
ZNChqyqdbbtX2XEGvAb2qA/ea0HeT0ywNcyw6a4B3W98txXnCz+JnYGS7oF1nN/5MJQK+khKxX1N
ie+v3IRq2gd2hMumfTWXzLtE9DTvSxbUN/NrLzrxqLKdE3CvYK9Q4lknJPwd8t/hEX3pTHA75cXZ
ZSV/ODb/SJm3ivqJ+XUlpZIT4Poa4+Lf6SUhl2twcNZpR49q/guKJeCuklOP84D12S1Jsatl0cSh
QNiWGOTyEJiXklUqSqra7Jx9oApRf1/bhbzsvj/Y/SobrEPJo+2/ACxsGdWFnxntyjSC6ThOEgeR
Y9xnhoIyvIHfKKiteWHI+lMVXXDeiJN2PAicjLspijhJcX1EBUtPkulYeehc+AVCqIaj5hcJK0wz
5AdD3AQcpX2Q/qFl+2+IDuY7Zxx1KkXSucMCudDATl7ORphdX1Rh4nEurb2rchHSBozE1oiZ0C3Z
MKMxhN51Y8qtVq4q73yAbnK1uDZzb1rydh3G0nabAiWFJqd3NXyzazINNitT0veJJUMHdjo5+fpA
ZpAk1MPK8YMwRXK9hOjxEhcfiUyNlH/04CzIeKxfAI5oeHWijklW+k4a4U6YydznRbf9ch7xaVJC
j/4PS0+NhzSSbMeEkHgQMWU3diE3cnIJILP1NZijk1sjBLNQwJgKoDhONz19heZd2p1G0yzrewIO
Q8TWZbQWLYrY+rdeTXozr4RLogoLuTaCXVqeVE3tI9BcAN0ds0kkySgmRCFSm0X2BEl6rdOjVuOM
OzseTotEzG8ZPeQ1foO6TRW1JozWbA8truibUBqAvpLgjxwOPuQxaqN7iO1djvN3eDmS8H1W0cdx
aUdHeSTXnBwgUf6l92rLGMYOpPkPMJXkXIdSAOXOiZDFKGZrBEq6EmySVzXLAXCIKXvPuZbZUC8b
/PuGeuQdDqBN3isHT/O3Pv2iou7TS5XcwUPvKo5STifSM7NMGEcYj+91jOQ5nwKRNNo1zhzVchN1
Wlrs+ibgusjU7b7qfr/p7UrrcD54l/un96SfJcL7XDhg4XEr5NdikhjEu6QxQsj7sGGPNJJ52xXq
KiriqSE5qBy4JO+MvzrVtDribbRJrs48/52K0rNXep6yBbZogmPQG4sN74tB1+/ADnBuHHhQUSe6
8TXs+EvPEmxq2Kw470HattsqpZh9btE1HPwX/7ApudvDqC/2QHdA6jh8mPgtB9IX6PS6aLMcz891
B4YMUeAftTuT/iOFNwPxvvjlSjJv+5/wss5JmcpLia4aorQYrxufPhi7VtobLhOs6e82jhEv7MnF
trp0m9fcen2VgahZFy1vmH1m9WO733PN0PgKH+WbJxdUDi3PWlmQ6XDCurlUL61EGKOLKuCZJ0St
z+c/5v56xcf3w3S5qvnFEyTDrFWcTwQ3AeRklyP/uoXe8Dkonq6PkdKv3ZshKCr+YzajM+EB3iks
hBZEjkMCpaOSTuBxs6s+yZwtwePn9FOa0tFrj4Az8Zp4mjjmWdofVE3hUJNtJ15t3gM65lF17EfH
DXk8SDGKZw8pwOJ7ZYARb60nh0BjyaYVPql13+bakp2QD3t01JfGLjXvn4hjfOCo84OgnLFhrSLc
hVMZaburb2rpz3B/lTsR5tSiu5lDd/1iedZBrsgls/1g3SrqwQ6ylSq4FMPh3vavmN+eV1UX5dRe
Je7Rhu77weJkYfDp7JJbV4kPlFTIJiVEmSTXBHeO0P49jk0/hFv+b45qQirmTn9sTseWJjsc1CNq
1xfp3x4mrllABr52APNWrQV3d62kAgJ0Jgx6OladNg3A5CGaiE8S6KfuA1vyP/kKoOMHhGzntcLm
7NzmPLGw+d7KQPTv2tojh5z57/40rDg4MwcY5fVFkksB9phOSXcke3BRa5uliJr5GNRiDbjY/7OX
AV49AeP0e7kWmwmSx8EhrbrrIYdzClLu5+3rO4l7DRf6DnyjYnsYN8eVXcsnb5GaZOXcng6OGkbA
ZbSWcJtVp3b2HjtTnVFh8nSDJ3cowU//L54TRx9uyvBYzzLldfvw4WBBXD9Gli7URI2joseuTPLV
eFpCP4R5gOheteZcp/1nyvhyyGWiZ35HF7W0tS+UMLB0zE2tLe42IZ2b7sJeSIni5B37x/WQxBVO
hJiAFug0QDWfHzmeJDd3XLd7BGqEjeYz3Qs8nUIp93loBsiSRO0Z5G/yzeghJINtiU72Fyse4+fH
EcaRh79ZMOL2I+ZSzLg9g/jgmvKi06N7gX/qvAtuW/a8IvNNPf1Sj3n2NT82v9R4VxJ4pvxfRGid
IILhgMlGP96lR+uQNQ0Z7KEMjEeINbbiOBhxOK7ACSlvAmH+mfS1XyitZZ4lAVCjEDrORUHW5xp2
TFS1OgPytrVcYKmDrHtMnXdLoLgI5AeTdXPlq4voNfoyBRsOmkK+vH+mb/eKUeExfwfSw20B40y8
tX3W4OuEXfq35F3ZI0DfLMYqfiQcfC4hvPTLSS2M1bD0q4qCBKJLV1nPQG8jF7/CokcnDye6ZNtk
U7OufwPKeXVN/q3Tw8Lh1BgEyQnLc9DTufu2VwHmox2sweAuSfIQ7/hEDrg1EpVOFfQNDmo5J4h5
UDmbl1V0kSmrhd27DaNB+dZ7c6l3SBp+V+LvDuQnpwBTEqnIH6QrEARhP+prPH5PQmcbqb3UPYEC
ujLh8WiGiTu6jHmFOMoDDA3QdFA2pm+xpXNu2jBhoOtxA4qDtDKa4zvPCXQwscqZpcvLooiEKyp/
aWcWOcNRmSqYnEWSmgwEis2Xjlo4BRjNaA2AX4/jps6nlOKxBEB45ftJTexafMDhSgC9GyHzoAIZ
liXAC08FLfb5K70ObfscbpcMCB0Yv0/35f6r7SZehlS36+uA8BWQ9sfm6Q6rMmf7m/XJvBmItKET
bwh77Xm6Rf2jWje1HS8dRAXrkMR8AgfEEe/IzdeQPbYaW5ghAKH1ifq6eI1zrsoS2b4e6fKugv3s
VgjUV4I55S7UDfPhlUs4CNwpYUTnanptfdnuPGlYFiJGlcGHDZ3oZnYNSEqE5eKlRryUPt+zLjtc
ZM/lPcFMEfWItcwAnyNgybKGZBORO0VC3AtE6EFJAB9pSMTZzO9dJTNoxDZey8e6r0AK5kuBqiwc
TBiWZOd2VWs3Wp++spd1cQmfPnqFVfEk1CGgcyj68pDqIqIFIN0p7m8zLS5Jz6Li3Zb1jTU3Ck1N
rcfg8iSWdFKdewFUYiZ8fu6RoZ5KOHKI4GO+nSR69IQOLsRpK3VbqrMMw/flah8iabg9ShoAplvq
AgnIdAlSFsR9u9ekFcVcZhZslSJ4jMHGsaJbowKQObT7eX3etN0VAkl8H24s36kUTn1WdP7u6FXt
IIrpQMDuzVqaVPMVMeyY+P9fIQH3eXixy4rCU8JmtT4qI3vUHurjc9k4VMElkGzTytDpO1Lx6mr5
MeEJnlymwBdptASoFjf4jewQGCNtoOAElXW6j07oDk/sbUatYO7/B0B7BmXj51FI1p62xthbf4gH
V6C4+TsOHxhv66c2lJC4NicGjDxE6nvpKBdRwSZnLHCy1ohgECViHjE6GEtupdeDJfXX+1sD1TbQ
ibzHBi54SZ68PW3Bhmx9aeeASgn7Ed/d5x9VBEqwYB+/GpqzNBgR4nAP/LO2yQZkjBGSt+6f8EZo
lpFhBVzzW3NT6jhqkEFWfkwE6S4fFAdgnqNbzm+FHxfMwLBl1XHMlyXFf4aCusjBg+kPBy1Hd7S6
OUzLLev957ccl/BjzschnCo5Rs8aZIevgH3ZrSDcGqQHyExx/YDNqPLcrskqB3tqHev7aUKqOhnQ
0hHIE22H19tt8N4P/so+aZatFkjKrLCchUjumHwSw6j3C50Z9iQh2qckVVoZK6DURm6zV2DnAGDZ
ak82Lsp9qex3GFMrbMHSPuHX6wkbxOrEH8vLAnzWgE97dvkiXmTBezDgpmiTYjd+DQ0ASHpyx6uT
BHYwsFUiuoMQQwIkCaovvSAXCP40uNHJ3k2jDGdZDi4eSZ40XouwSxWhi2lVhXx5zs0bG49no0XU
lRB/RPPQfjcdGnhdNxUpg70PaKXb3Bew/oaW6BoSDZja+5NwujRZ4XRmrDngA/Eb1GkZOwb0yr5a
VIUUUEYbq8XINBLlp3g2uBcAq4qD+x6KIrgq50Lxsny4wCylhCh3F6uUiXSHBmy+gqCL2dI3trnq
DXI7WrJ/pWJCHmH0Y+9271fxB8n/M+2YFY62wcCCnoyYPb/hVLRFyeAa2sVcCwKHgLaC+yqszK84
lDs37j/6TA5ZwlOsN8k85w+GuodhMGFWS8J225ccPRH/3DFOtgpvXBciaIezzy8fdM/SK7TZZRfI
4LQo0RZ6Uscl8tEcT7GAuXL42bOw8d4O5aOAvGJjLd7qemZAuAAOaVAkPU1DDI6oeOE7xlFWhYiC
31QjMW5Iby0rWm4oKi8Eqm3XCR/a8hLvVfjdM0SKF8AJgZf96N/O1/Sl8SzrdQkTM/jq1w+3Ts6Y
1TF+QESPRGD6qrTzdd9QajJ9t+jPd/QA7yOGNle8MblumF/Fm98gynI6lyxEZK5wSI70X2Oh71LA
aowapF3diIs18pcHaIgg8RfolfBv4Qpqjd0uO8L4B3o0cjMkcB3ofZOLUxLZTZ8oE2kukuShTUDT
Rr02Rf0M6NfI5iRhQ1QoDznjtjy5sse1koZl3WSLyGasZBKNTGNLYlUyITC46lkIKzbjW52zIWle
KzvFnDFVkydojmFwniIxqyENkcZtOofQpXhHObj7DceJuUB8N90J84fkQQlIAsfTlkLHa6hOA3uV
yAHNizM0Vkw7EjpX7yhjM563LzBpGqac0IEbyhKNbUxnJ8DxHUYeJ6+7YZy4gbzeNgRJx7bOCIxB
2rG49XNxlUbPJHPi+4WXRRz7sf3SRBAClDH1pQHcAJRwuyFn9qVj1vMV6ZF1MsPlA9TIZifeiFZw
nTGAb5bc/VefiT3dcCXIrAKhjjSxwpWHwcKeDiDciIX7qSWSC+39WzsLmdVNOvCRA6Bi/oIjmgnO
TcUgYSamoKnRXQLqK5H/PepxFqjuZl+p9oXp9P9IBAus7srgKldKVUPWo7wqa/ruB7xMxg+Hi5Yg
sMBXBEEI01nF0k/oWqtU//HsoxqK8MIN5XMESGzFhbVPYapOkRaIVVB7iiSlUEqM62kOehZXf+oC
dPI1wRjhBDwscIaSTdzovSFKBHHppG+Y6A0vRSmasaQAtE/TkzaTIe64GZkf3GaQ1JIC6Txt+fFK
ob41aECBcpmYHIbatVFw2XcBz3SK5azcbGSH8FnRaxT++PPCtrbc1JqN29Loz1MdAzHlSmvUH53q
g8Xsf8oVNmms5xXtpyCFjJb2v6EwYq3Ztt5EysrsB4EBm39TQtR48mRVKkNlWpLuqG2cMl8hDrTv
/hkxu0cL0tEP9Vdi/7xhV1XQRI2EY1a/XaL5PPdS6LFhVJ5cp3iuQzVv8MVZQLJFHfqaxM+igbg7
iuWF9k27+OUErCV1ipLsqRAaM4FLKlB3XKICuevpiaQjzIsvEdyG91YnlkdihUJ24qkLzF7Q5Mxd
CBihNW6MLt4dHF1jiwNIRdyDNR+zXs3sEuo6tR4NPJuzKGPAoAkCN00bpf3MBQ9ipTgOGqtkwjvN
kSpIb7uqjg0X9Ctf2doRzQKsNVEJrTwY0DtLZrpDO6gVJunDo9N2OYDAtl512taTfmff2qQ05m/2
gb/ZUEFbs+quQ05CzFzZKj+/dt2Tl9TCoE8wYxs5EmVWsK3GOoujqK7/8t8+fbtjtW5JvWbRfe3Z
mVjPFTO7XEjUw+/1MY31wLKpGK3B9xq4biDIQQGVeQds8c3y6F1hZS5MvpPHmMil/Dp2TN4EPnQR
5Doaw/HtQ76zxi4oJU3/PCv5dTMLCnqOaVJCI9J3y2fykevv8uscab0W/WxgNBbVzx54irgtnWBa
44ljW47u7yzmmtMXihram/xOIMOF8pso4jfVVVeAIlyY/39AODBUbgcFiLdmFmAmN7v84PeJpl9b
IqMJ8JzO40BjYgVvXCJ5M4z3hbWGzamcMw7jSKQOp6dXp+oKunsJuR7OTSG5Nld4xn2fijfSTQjL
RADhLfGe7TUWhNl7ou9mxR7/kAv4AMhilMSreRaZmiQleN5csUgJHOoA4NfsNBijPT4PfNfjoPKH
WQ8vwIEuq+TlkQ2usWPPpC24Rk1IhxQaa48PG5judI0n2ZIFEInsc6quKjqEP4Hw6OKYutKQmRx0
Y0eQZ4i9vsIz2bPlSAUg92VrfQEBKLqJKHxzcnqaeKFsvcgDoJLLj7Oxrv7/BgqHEeU7WtvHMMu9
Goe92pMP6vOuYPl8mQzpQPBafaNLTCFRsHQywygdnESlFNYXJpmnq5rzv82lxLLigJPmuWJyH74B
cxcEpfhhnjmLI361INHbOfi13dL9jWNzg/q7V1n1iBMnnTOWFu0AU2pppdp/O6kcbXgy/DLc/kgw
srD4f4LdMrQAmLXOkpQUWMUnIrIwj6gxxG6fb3nL17k50tu2hn/62kNhJjT68WAHKgQkOGrXltdF
2uYHxyhd3WY3C5fiprW5DSrpZdn/Ob8GnAYLaeb5h7i0Q3CfW0/KaCj3V59ACoN6RLj0sJ8inNCm
sMGW4ujg+LpfxRfBTuJB9o2GksdEhzcazAoIliTEbiciUc0jVraR9ArPSVy76j/WSGxxw0ilSoyU
2HLEgwV7F/9noCjBlMvIuUe+m4OJHAgKeGNHrQDl/qeUIT62EGtqcqkhRsdPCnYlBK/LdQdUMro8
8r1iEk1hRQO20PGHhZ/SQABlAdJstFavrfRxt35i/Z4XWqNlNB7j1z41e31sU94FhcetFvgOG6FP
lCbaB9gUFyx9l8GVqoQ04zo4QpwMq47/vH33VqfsJfy8OgTk52yK3YchokAST7+xCbubZEWUhw3+
d84E29MZ8Nr+aQoMDpvpt2t8/oVKfgDAkzsKGveDUTkhA6BA4flKP5CnO1kW6p/039t/3AHFCEPg
duE3L8tY7mi2u4AhzGvdj0R0zLr0B782a/xm+UU9drndhvzys2fANDuf9WGvFz2XkRjWwcxknJ1L
q93OUhLhhYt4oRjWpGR4AAtV6iL500TwfnRcu1Mwgt1jftx1H2cb3elyJ+e2Nf2CRvbZqcj/g+ko
g+oeQJabesY+LkKbet+HDVPpw2Js6/ffhe4MyrlCpZ0FTAeJknm4dd4uW3o4s4drD/PvQqhwL2Uo
0t0n+rVqFinmsbL9WDYEgBZ4UFjWbKX3gFJDgsVfSGbuCIFZYY1DxHZVQU0xupkv13Nt4nUU2NfU
JPce+xYAFBuKUnvXBArd4gWbzsu9vJ4VN+yDZxAIPR76luLnSeLhpZhbuSbXAXyDRl4vbrOil+O2
RWvoOU53vl7Sr25bPRmY88L+A+Wi0wT+FCPT8R0zCH5yyEhrRkOeUSuEzwuiGzozftL2rWbbQMft
CRS/FSqFwm4cYcx9TVfD6jlS5fjs1wlqScmE4l2RsQw7W5aCiKiI2+SooqxkjFAcpv32qR31+r7k
kJm3FcQLDXFfh9djACHoXDeUfQWAYBx7wKpWRoOsfSyRUgUCWZ4yRGqq89ZJCOGKsydsxlXHWCzu
FtPZPrDAzHm7/HvWBK/B3Hjp1M8VJUEnBAB6QjO+vIyyFBCyw8oHh22ywCFwB4HGMRC42AKDvX7I
XhoAhcoewR6E0DAJd4aiDbgHTDIg3w8/VqJ1jpRy+Ia54GPzAnNA3+05bqTG8UZroe8bvZbU8Xwr
c9koVzM20G2BcSe81tFRBglX2sp3BODozqSxksw8ch5ePWNPYGUoPXcP3WsjmYoXeLG+LYmRxv4n
TDXOOCb7BqfDbA+y9dgn4EYAprMY+IujPHGPPVDjuUEFLCP5KV6qQ4thLjcJq0EnHGbf5/7zU80d
RY94Ol1fBEVlBYLRkVPr9G/qwxVSDzCLbrnLPI+1T8q8zX1K1SnVXNErAmN8Kn8+ooFMcjMkPwhN
qYuE6UHOYrE5ox4VGD6Rf0FoqgbRcKfkVo8ttRQKTR0d3y8nGLfgG8upDzNS/XSSfiVhRT4SClye
z+PKbpiDvdvPMGY3FnP06Lhgkk1Az/v6JrYHCJ8IByWVnQOVcsmMG8rIPq6e+BbIm/VIjzvZn8CC
sGzIYNIbsEx/lkIks2Y39cAs5Pv6cPCdN4zMUbxZyH3gTEdvyzljexvteFqiPMn9L9vV53/89bWX
bMzqFupMLpdIvPjs3rXf7NYEolEmMM4mUfZPSOWZqkSp9z0MOH2MA92a6UD5EOUbHzUxGp/ze/Rq
hr9zNnDKvGwL141oDLYa8P2SaiXgB1CLwRfm34ffvyvID8I7TxTNkyc3IY9z81L9RENwnZvy3fR/
rCk0FlEb6uDPDD98U3fIzc7gnIR1ZEbHGYgBK1SUdMAfA5o7JyPYdsa9Cpbc2nLDRAADcZR6MI5+
ZT0oK88Nunn3MiJZNU3ydZ6SVypWWJFhflECQbBtLxvtwnsp1nZ0r1WHgGEtxvYlgIXCD7z6+YIV
PYxzt8HSb+3V6VH4AZp/oq+0WpqN/PdxZcI6acAaJdrhmStu8Ja6auWk7jTQyKpWeietXc3rHRWF
Rk1Mktk+4bKOvuvXpJujeMVXbnLbO4JvWqr8EwEWpU9eB+PankGuqATkcLrdIAnMqdTGlDLJ7YTZ
DDT/5c/jDrlpBd2dbtVrbGQekc66ubXp375FNvmee/VvMd+VAO6zImObEROWNPiUq9FJ1rdB9BQs
so8AwgqcFvK0XOn1wCKCL0i/a9HWsMvoVZvqZ50XTj8v+A6MYHcjyiyA0F/gfsnWzMiAcKwy2NYU
22b9AdTaV8ghcu3fsMVvoJcYMeG9BwqRmmWMsiXnRx+BX8YraY7W5EXV8V6C/XxIFV76jVVwh+A7
q94MpQt19ehqivNsJKjB4XAtCvVrxkrFB6wFflkQb2LM0bGfeJNULxdF8ooC4mSDHnAWf0aZkPAh
lO8R7V09J0jS3axkjFwOY2QNys1JdQLz066/R+uojRTZavGeX5Ma29K9F0JZhLrk1rJYWNMVyWnJ
aMXihHyzdCO4OzE0OWq3Yy4Q5LTAjwe1uS4+4G3tyufzjd7He3a3nxx5MldmAqECj01spU/p38+i
+cFx5u4IFCuaE9i3CqYy3d2sz916vKwoprvas1eS5avCfn9t794T+HYHsfFr9iZdUlgWfZ0QrqSZ
ryozgP26lvu5BR2+6tOZyJyk+UD+ELafd4fI2dVEgRx0GC8DPCDRQgKSGBOSNMbG3WQplDCaJEzC
sjD4SE2wS9mmzF2o3h0SQJpy5NA9clpEuJI/do52eSP7wWBzByt92TRpvqjeWvnd+NvihW4M1v/q
ZZElrgkAmFiQpc0woH8xviG7R9lPfAlgxr1iA+Ch4pY9IPmx19vD0rCY/KcStNHvGlJIoDVF56Ba
87f5oJ8Q+OnnBmY8R7WwWIkuNr/Y5BiWP2i/lHA9hP4kF8qvy+CKo+WZaZKyyaPwrgu2eJ2X5ijz
VZZtUVMXXJ49tuzzh8bMvXOprfFsG77jMAUiufZdiZ38mwMqEdkQA1lOEGb6RcXdMK9ATICQUePQ
6YFjsteZeMQ17C3coKjUloL1VxBjhwRhce4WNmBvqZ3J3nKyHtaIBisGQWKJBkkOoe0vDEXjp4s9
Wzlccg0e4iboAdxvSw23UY562wvWPi63fW+6LM1Gp7iCKfZB6flAla4Z5fEb5m4R5bpUg97BC4ev
khyk/c86/BLtVM55IVuoJKbMBRkH9LygtntZxV8LcutBQgX7IVXoYajv8V3JMxs6PD+ORIL7+NMa
sBOYVQobazrMcwEjwuQ6I3EHec6D3+RMAwDCsMF+QhmsU6UrkeNH9qGDTkhb5K2IbzaRkkMd0Gmv
4hpGK0d81IN2AdKEobqdYZvRxWtDCKmklkQ9LnTwtDR/hzlIISJZXGJaFpjF5QM7A1dwF5dUDeVY
Je9/ukcugXJs86aYeVYVFMNZb3iJsTAbtPJur6yuzPPtw9512PQUsDinz8aYIvdYWiOMvEUbUWXh
lVFD7LvupPCwl0eiSXcxlCaD3Okcg3J0hKvCVdHXE3zpIGGZ2Zqi3KmQCmipX06+fLGsgXqJTZhR
Rc4Ix/zPzgef9ji0gJW0tuUBa5xnF/SyJ2C8WCSEHHDbQ1GCPUKIty2lOBN97LsgVuS8YWwSmOk4
fvva5/acmzyFUxM7lfPCoXP4DqnBei6jDkDR0Rhkf/qrMYHOnRpimQrAPDPQoSQrLy543GUTLByt
3GDYRmlVBEDmehADVYiJQNLmHLdGYIM6AcpYuzKFJA1OMiWPfrIZpKdrv8Eusox+Kvwk7mMlS+qG
fhiDiWSuxzbzY1lS8tky2rczKR0DPB6Jo8j6mo993HP2xMoNfSYz62hMyaH9JvbwChbuELsZVxX4
N8TPsxlpN7mWjOnNTdNk8/4NOrEM9vuqPn+eUWbRqcfsiTAtS9T3FLy6HNnWJj0C7HzOHeP8CGfB
WovYM9jZjEjWQmUeHryJUJuhaFoY0Ya2oMeerOCTFxmpuipyjbWAbSj+lvQxOxFnq4e8DKYlh5WK
4BSws4CmvUqYpkl1kHr/2dHBIjv/R8VH2V+HfznIb9XfepDgXCdPib2YFaAchT56wQ4cO7t2fIF6
lEBhBy1TK3sfATOaCa7rjB0UmdZgPCRlo+zPdAo/fXB+VLzBMx1Ui+kOfEqqH/ldadSTXcM2yEGW
my1YBlWiEEAcs8tj+Mzi403obNFknbLRYBpP61xB1sFEFlbc/+MHJ+26KjcigVacLhGOLNNUYKwT
LM8z5XvWfE1KHmZOsuk8gdQeYEa4U+8oXPAd6PcDN3CYsFICGCu7BVYmDQfPjzk7nPSPZbvbXXaQ
chn7+WMBiXa0s/ak7dHmNWKLOF6ung+JIb+soX2VH5AitYoU60PfVEJYL53ZybQmY5KSKkM7txFz
D3hmu/C0ooMPm+66FtHS32tvQmGVlu27xpPE/PnI14oWEmEtuXNSgY2BZohfnS9lY0l56Rxm5qSk
UU13335OTyerULp546T7vfP4QK6Sa+MDGgAjyGD4Yaoq/HdZJXbwpshJdKaYJ4J0K3uB8RML5ywg
luwXeVe1SrFWZLJqf00bdsfVWAGXaUsxWYTTRJELjddiXoIodnr1SJTWF1+5UFODggNDVyfVJn1X
yDXl/BMDLwbgiddfrN3l0cMV64gulvJvdp0UC0RtCQnVPgYOV10hxvz4plAMKBqV2zq1Zwtf49cO
JFvMhIajaGTjaoEs78LUW4XBY0gtkUocHaj65CUwJNN1lxdo0lxfINwVSVp9ieH3qdNrLc7Cuw0K
emNuo3UgLRtnVJQNgwpv1am0avYM99Q7z+HLKQ6U08257uY4Q4yHO+UHAyIf5wB6JDFKKtnO0kQw
iDTYpo/odopzARiEY7YGJc5oKFeKn7P0pXiNK0YzknWbkCrym9FhJnNxmZwzqvmVIoO3Fu6wLGGj
SXAjcu/lRKdFZeea+RbD6nsQlrWcuG2QSvQVDqthwDBBXc63NNHAx+ESH+g70+zkCaL3byi5ZWR1
gj/XhlI7jjmxPY0AFhJry/LCjoIK3rbxkjdBCsd6f33qJqQlmJfnrliyz8U9bPL41mm5e8mmUH38
x1vSNHy9szeVHiMxiJ3eOqJPHDbw2XZ+LXkQGtMV33xSDGj3jqWhkeL3hHzsf5uuXW5boRBwjPxx
BlSPILG+C1prwus7QTUtORXSPFScg+aFnPjjU1o808xoHtyhqGszscD0BfjE/0bDwDmJs6u0X1ye
yVrASFcJutRHj+pxY1aMLx1Qu1gOtWpRepTPa1VtPsoXz4wHewFlG7USnJ1nN1oDRsba/yxlysjk
d9hOuMcHE1rzA/yVt2DYDN1yjA9JtVqRwLUY/9evYT+LBLPbS04YHCmIc80xXeR9H8JKFr49QXLn
Nxow/FKqyQzybM4Jq+C+cH/iDWe6aURn7fAAbajyF44cxHOzknjgmvkWht3fHw+j4suR9KWQlGze
SSMFr1MOjelHGNzDyNcgAT8QzGHKni7wIWe+pT6il53wIoXRs5mX551CohpA05SP2WsUAR9o3eiE
YyGSNqO3y8q6Q3MeXS0nrVArbTmOldD1z2Qh2KTigQz9gby1NX4doWE3G6jLbtONDflfL/etdGPD
JVHEVxn6U8+Xl7rKUrHLi2LjPCaPow16DzLyevp3wBLQXg+x4G8aWmPyGADRIYQCbS2LYyrH6ssi
qzcIc5xrvl4DbEgHO8rVsRbmFSIJe7h83y4hKkFfS1Ezql9hVEQ6Myz3KZcZ5lWw0B+9h/2hhzdR
T1W4AoMsKnliY+nc6190Ttyj83KyZrxD/H/ZlNQekbffjCtE6MzzZBd0kdJ2GZASnRXozLEAAXRt
tu8SHkV6lLbB0PrMx+rvGOyeObT9wYk1pL2FeMQbVewiHuOsRF2Fc73cF4FB4n39O/Ku+3GHUvFd
bAIf/UQittIPuigynHkO2uFMaZrL/OVxva8D6bIcY+Vqavx9x+Zw0VNPMT76BAz3pxCWMNU14mtZ
IiBwv4EhCjgjgg4Z9VIkleL0UtRRW+GrvHdD38gShjp71WkhKsfFJYkEF8rLAatMou4gBOKXjm0q
9Slsdt1tJa2a6sV1Fl/ktfpHsfDQmMkSkEPKRd2msMi2qGSCVkU8v3zFQnpdUupoNkzGVH2ctHkK
p5BqODdohQyR8xD4frPyOmn/2qX7uNnaGZQvVu7I8q7iGYKSRrRPv2tS1xOgLXRcvZddECKQIfl8
x7rZVmzAwmqkCJgGoWvViZnU1mraN3P93wHqEJ/WAdJ/KuwJ4YmAaQrnS3TPzzfHYdrnYTSWw2CA
+6eAmFeZeiK1rsn2Mkl6LWxMlbi+ZtIbPpCptwtWCsf9ZnX1ftKVjNEvaw6z1UIHzMSPdTFVf4mr
4hj82MGCeMOg40XKsspaIWt3WtL9Lgr/KU75MeNEXlxZZ3PAmrNFGkGF9cSv/YMgqGN/Rrc8VrRC
6+hhywMfOZdbEQffi1+CwTvgI2yZhJrBbnDahgpsAq/wR71dx7bGLffizI8c2OrcG41ibvSlpdHT
qr9GeIqKFiK526FY3WjGIoUwJdSCu7CUjVYXDA3OstxRJE03SukTrcTPSxzXDY0aJLdLfBnjpb8z
tGzCNGh8o+G+Tis/Z0dpPUjB6FqcuH5PagWBDgIxTXn92/YXU1NtbKl9NJl3O0qQWwmC1M+51ttI
jvqKMk4pxeupvRKpAPZFnBprIbCUoLrxn1OSA5TBwcHQXbb8STtiC2oAnnHg4ikUPDbux08ndI3z
dSKPanM211ogStt4ii+qxcbLIAHjA7JrCpTeF41DCvxtWtYeMmYx5XF3CGiJUn2VgoAf5EaPtluQ
hfIQtFUr9vC0IG9QYSN3gCZuUKkmaaVq/vvzJ4rUHSZlIs3+iUVw5HTZBYfZRXhRy8ViI326lm+N
dPa98BqWtzo9/LLWTmj+rQqmHnvuG8DznG3TNRV3QYD1paGYRUjepSLrOS2RaWJEUtPAbWfwf6hr
z790g/Uf8bbo+QFBK005CVN54GzTsPHQQcen/v2M8OiAV2Qi3dQZM4DSoNBCYc5Ry8hD3XjzETHw
wiR9BR5tKKqPZNUXj3RjG8pZlkbh4oXfXCs07sa9PHXF07hfAZBycanr3qRXOvUbvXekwoyiWpwz
yTtHQvSKjP5dtD1Fn2t/YC5DJe6NrOY0hDXKZpf6VNfmLHaBDJQrueKe1SFF9yHcKAiYXGUhkmG3
7A++EEi5fig785hXdyPuqXsm1TNx1sJMJbp4/KWNW4E+4v1YqcaKBSThlTmCFpgWGpblDbt0JdfN
r+S6eKzlsyW5XwPwx5yH3KsLr1dBmAyw5ytx/qT9vywPeBxKtNN7srksRmdvMNmfv6nloDTYFQ5P
bwjnZBWiTKBjWGTlpJPllgp3Jnso57QzIm38+YGvS/OVKSZT/+gJOzL/Wpoes48lnE4voROylJK8
XKOkobkHdnV8M9dJD+vP5a1t1/gBfQTXUyckOhv60WkPFvMLxzuyS2JFSzajdKtkX11A0eytrWtx
BAvyr0aISmMkgU+UswN7d0467iHPMGlR5sXwMp6i474Dhn5bgOYp3JDmhAM+Xdo4yvr1jBWrlfCE
/PTrqSMsi4sSSfC8QJYddMq7tJ7ucd/25eDZZEo4RWDHJTdI7uL5JrQtzI2aofWdNMF3AxwYR9wD
qdJqEw5Mu8FoothZj6GVGPBFMIXXc8GgWKxz8hcy99z0NKp0HyyjmWzcJgExGm83jZ7poUZQCYj2
XiNfwNOcM31mChjcg0wXSPuYNE35NNIP6an1zWfSVO3a+JoiUrYNDOC405+O4dJ5WmE2AR3RCkv9
DVndPFQG7jTSqNb5dPTf1cl5f90G25Dh3FtjO9W7xXz/LBrRjuUTy4ZEvlPCR9MrfpDPENjo4vSP
REch1RnvBnp8TVod2y11JC+SeXEQR9cuD1yskIZ2Fzf5O5sTMvmyWSg6++IjsERkRuJRZw0ppTas
mRbO4gLKdjlEpcgfm1pZCuNVi8zGXGnkTDZG1CDqW7eSVq2VK57KikDcIOqXIDzDLiX6dn20JNqT
cKXGyYGdvcWYVppTjksq8j2vvBFcMjgpSW3MFcYBWpgjiWKZKaNAmWMB672/tAAAOhGM4jKHWYoB
gfgzQXbCkxhoey0zjogjzqb4loCWLW/d6D28ZPXn7Miz9pFtaFFa42IM5Y2wY4iO/GYEpZwSUrJq
f5wxCFS70zV0JqmT0o8LGPCJaOf23oVtelArkHRt7j92o67ev3+ccV9OeprlCsVjfWVJ/gUSu9go
/WZod0RjSh6tHrCRj2kLkYU2cnNd+ZK8BWA5Qyw4oz5KQtKssXZfHn4xeN+4hmAJ6WEmYpvffhiT
ysVJkEPDJif42K2gAGLC7hyo9xfwxTnVo638jiSyUZRkk4clTcU3euaFWBwlqf10zD9Hfwz78dng
fMG9LZEUD7CEzy8JVyqhxRC1pv8BLUorocJKtWnXVaFAItAs7Rpq0SmP9Hp31qq5AfOnt8yqwUVW
ZXBbubYnolS6/ydP8Tevcpc/eeqbIX5blbYyX/rHwesEIUT8drqwb6PDDDAySYPaCaQjdUWbFMlt
KDBxiIQUSvYuwRrpbdzVTf9JcPoVzs+xx3S1RzEpyks6H9bLiNCmZ+2cw0lElNZF/zSOzrB9xbPR
vlixKgftCzrDTePh3tu+tipNEvWM+yRGL2e11wMleUDF2qhuyAqEStt/27wHRcA0mbiIXcvCWc+e
QFCJAUQEKF0lACb9MXWeBJXUZUOUSh9WG7L28XO/w76Af7XXYaHfo+ES34L4mKfEezl4yqQGMG5K
h3LmCJ+i98PsDOhDiyYXSGksxvfbk6YAY7nFP+h5iHvUYtdEtBx5Kp/ZbjNoOY6UXbnifLkzQtkv
S13Ci3JyVqoAYjPTWn60X2RyZ/DnHAQbZn40ASGEMeWRiWkT4P4Z0CcZ3YYa4fcfRmJNile+0VR1
ohDzh40YWs1Pb9udjvYSpy1kPuaPfWsgyBi84D+aw1xErgq49GBU+bapMaoLIZFdrlTu3fsmPKr5
LSvN2/eqL030K13aDJFq74qeIjnOaRaFq3fwkS+rVZ3C7iYQoSeSOMf1ju85pfc8hCWTufVsuy5/
uo86FuOmD7XdkKQV5s/JhSzo83a0pHx4pJFGk28VRxhVuRcUm1Mk0XiBkyhl0xfKnxJVDImrTzpP
QLXJL06Mqp1kckumXD0Z/cx2r528DCzxOZKHjA7QsGcz8fgHZsWm2INY+2F2VbHRqguuZe4o29lh
JivoEOwUsEP/HVyF1/IL/KnVf0K0Jal+qTtYmUbLZmWpNXvN89+l9Gu29QXm/ZUgmCli/3FqznzT
fXIrQDi5KMYztmgLVzZsXSkQDNfucsuVjwlp9qQProStgs4KxvQrGc/DCA/Pze8vYi90DJeStSQz
3kNVz5ZcHHrkCwxozdkZxm365AsoU1NlfbH1L2wlJmnNdn1rJTpikX8YVo0LQ18mtyrF91CU7Tt8
whtRptvawgQYx5aihVDrMsQ//RBNzfe1BFMCW8kOnMLB97pJIWkxIPd5qOtHnecy3Ans1aO9/ytR
6RHSaQ3pHIiibAXWvwBV+teeNf6Irk6xQKFW6HEiKOaiIeKDh+t/BfQrYhejYX28E7ewpxh19+in
pKljGFPFtOfQbhXQzhYoWEicnyeZlY0JwTQmsWtLxBOaVADO7rHLJA3QVLSstLpgn27eACxm5j/3
UdGr+miu2lEFowhmkrh7Oe5Bdxw3Od/3aiyKh8sbx6fUoXOmt7CH2KTNUPQhdbPiwtMShEJROChW
mCuNYK5iPg6OhQhTpeZU8DgeaQDwMA8PxYV9IrkazrEBOSwTH8uWSXRdABVKXCep2mobZQb3D24D
/KbCCju2BiJWjiga456WVT4D/9NWCWWhftsqm6Eq/cafE0OdKfYst+nMr7lI2t5HOl7rj7dZQXhQ
XGcciZKLwGz330spDsR242IvLDXe1hlXXJA4VOzyd7q/mPqjEXX1JTP4+Y2ZDywnzgVs7Z+0hIE/
iQB9EHqFa+lUw/i3YHgQnxvVgD6AZTIRw4Nj1OwxkRw304w0WmZkMWk0V6bfqj0BmLv6gWfIWMGa
uH0ihlYvp+wCq0eqFCdqD4mf6EgUIU6sCRJEsUaU+zqb/NkzRwOMN0J9ZftNnrFtWacW1OSg/gZQ
zJV8/ViRcpV9dCO40DiP7vQ795qWcbPz6tIVTeN2We7XuqUFUOiA0nsUU/Ke1YHvqFVzdwH60fnQ
oDb7puM97L1OjgyYVlv21CaKo9HT5HydyuEUciKFx0g/O2feLIy3gk3NOE212aTf5GHOAFj5lFCc
+LCEPHqldBkVSVY5nWlNsqHAEUtOH4TSptgsBUYLdPm0jFOiT3W8x86LjIoz2DxAQ5MeT+qvv2GU
mGLOcMeu76XUAL6B7SSrrMPbwiOP67aTbi1g5gd3pleDuXNmZX1Vym0FVJwxPUe8d727CYkXAWZO
E4srLDwAo7vK1pqBiloIbyEq3ube/O/D9gmtZfkd94rhfQe1uDYcNEGylRp15gs0A0GghG8RHkBF
npgFSyPjZ8rb1BpCbm0IiivQLjPlu8wUNc+oDioOFul8AeQFVSxWzoBwIvs2dyTY6ExwncttAPze
DTT6l0WDRwm1H511bVZ86xzHB4j7+NIONM7el8XO1oJnsjPBXC/fBc/9HzFnSQRX18+13KOg/GJh
abFqKEoGmsJa1fwsQcLIWYzpgmgXSvo2N1bUkY6oIeMPaAzsFxgjqhvMu8Pqhc3nSGylUOJUx0yL
WHtAaPo8HZUwdR/xELa1AXWMkfIIAsNCVYAMbptvDg4/Xmq4sQe3u+VqrNEBsKLQycZg32bCKeSp
UOJ3jfsLA/qttXgKf/u9Xty5c+Ay9H7evCBJO+/GyB5XPdKDi4sH8v0CyuFhmORgboHR824iy1Kv
H2Pakz4U9mrB/MYEHqjvVkYGoQBI4wEkVVuXfUz2Bm/TxpiTn2iu1pVHmBWmw2BPk7QtLLdlqpZ7
+OEe1i0m4KwXJzMKZZK0JqZcu8LzTTJJ0JLcxbMKtfc1+sDt4W0Y85WXiKGAl5SKBFJrnyTyIQFF
asMzcFVtaOP5uSJ5p1CkWLwLE9eXxmo/BrIP03mAsSVOiga9iCT9xUkOqqJujRnggWpBEqOThaug
V+mjNLak8X3Z34aXBBAADgyPOq2ZUOv05mIDpjL9Whaq8MK+f0Hkev0rPYugC4CR7Ih0onjNTHwM
8Zin0kqbBBYVc2BnM2IuTAZ7rolch7q5vAyeOfTsgu5meSlyldhdkT2YTmrZHmlBiwRyqGFP03mw
YNU6uwOtkFnbh5A7zmmOje9FXh5OnVLmreDqxpUabU3Wl8KGjuN0m8pw2OQGe8+ql0Dx+xbVJNM2
Z2GbHjjTe234f1VdU5jneK/GE2q3KP/6MzUI1i2AYRgsWDiA4IOlPeia6xUV2lCC7XsVhu9mpvD6
eCTttEBd2FHyOFhTY8hqdWn5d0vht0zO78gUeN8FaCLmBn6ZQo3vUAVMdh2H1zXdLieW3rUjS+5r
IXu+E/Zi0bMHnyZ7LalY/sEf6J9Rzqr08R0yk0ZPvPXrha6Oj3vgvkd8YO5eB/91sZBsxy1AGSco
WXokGphzfJocEbqI2J3uwXoZlNjzbr3V943G2meBQAEsoVa8XNROir0JsV6um6s1UiAlbnI5SqL6
3mHKHfLgWOonEcqEaDSLOLTjL4kEfBZlVU7iDj2kVu2K0rpYYScynnPPkH61QRDBAD4ERpAM4ul1
Mii3GAZRDmGYd5GS7Mdu0Nhjwdbyd3sB82FvSox2Uxvex+nVFoBjPqBBdEbym60wSjIFA9Yknlxp
Q+PAL9V8RnOwzVeIcxjCMIJYTCtKFQFrU8P+yCDVGQqYAjlp66+fU7upjYbkrt5Flhf+BVHEcDvC
6OubzkcqeiKT8kD8L+D3SEDOY6ilbfOnVXx4MAhIGMrm3mLVJNlXCSNiWn4uRSh7EFpUgdNr3VXC
CktyJ5JJLP0QqLLuzpmxA03iZK1j7bJ3pcl9iGl3QQMMnBA0TPlWvStgna0iNdd3d5Og4+HPJpv6
enNVTTb8OGC1Jl5lBiM3mOy8eoabVpT4MIcy9p+NT+2uPcOytd5sfHY3kmq+hcatKha6UAEaOhXN
YUCQgywRWLM+6V9cyLaZDwn19NwN8OT1AURAH7nNkLgmbWa5HxmHKL9IqrGZfHR7l7V7tLADZW2h
et6zmHhgSF13GQFWp0UAuJvRnwG5JvKbRinDPxhpp1OpgfY/9zdsLfBBYFaj0cSBG2jJuAGBUAoR
xXKsPM18D028z6cvFZ/vIEe/rVhDRNWHa13owiWtZEVNCTxqdsrraM2efXKbkb4ar7N3TsDIv/Bc
vItcjbojEV+mrQprhxcbvRp7kDwT6bIu0GT//HWqCEoVE0+yPFCVqzHnf8kzA1xe0SEJFkjZacp1
HFenKbA6ZXrLCJHUkhaiDjOJYQ9HvvAKVzAqe7IIduuhBxUOpDHmxrGXPOwqC4j13w9lC5On+Ni/
gf1W4q4235yFNegXgi4NAYv9pfLkgAbKsKLJNibxGvb9v/WcQWP2h0Mt6axpeJNwJeoSZ+ne9X4z
VuAg4JuxFk6oFTls8w1KraRdRLwOsd73k1bWQeAs+1Lmgm/zpy9p1tXtYFguRFWw5mQtpMkXqDKR
ctX+yyU7/io1IflsVN8lWegLh80KSYMSaeq4SlTenji2o3a5225P8i+MlEWeTyqdX7OnNqqDcAzi
0ZdbxCSiYk19n0Jg6p6oOi+DQNUV8b5eZoP2IoZXHU1yPFEWxKN6y7AW4HSiTc4U2mGFT9vuY6Zi
Dylyyi8L2lWdb7NkiyrThNEVKROr1bV3ObNzGuoMavm5pPyGKlQcOn10IfnsKI537PKS0wQOlQP3
jzhzC689gFCXvCY/RpLZC/aSRggdUfvzimrb25EjzPzi2PJhLXzuqjtZCbkGVU+0o7+Aaq2Bcea4
jaZCee+gDJ5iXKqYDbfw2O46Y3FhKhRULxdMCXFpX8hFuum5OgHqJBSCfdSHQNFhvJtfcLH7GRXc
N8rdllmhmqt3msGIaUI9udinZzo/SqMuTNxSTZcIev2PO6Dp0sWAX9scqEIEr3IUpyb4OK0z6Jv9
B1q2AbwnlhkFI+tGK4jOQdw19K1WhSB1qJ79aUVUi15eJzM59Y5NMoR3cu4bs00ScJxvEgKYdISF
MZ1Nzs+ZKiEABKLM8U/ARBxBU6Me8rLjBiPD4t0cX6KJ+lUaIHyptfv5g7CJqnO8sgZMl+OgTyp1
o7LhNqVtZ2J53LVkudroV872arq879PR3P2xozB1rqfMivxfewl+i+P9fd/pLxgJ6HhYoe2W+cNR
mv5uLwKyO8cf5LX8TRwL6QGdYt9RL41C8fMdVsy6UJ+qFupJs/F6Vydx26Dv61VDBnYr4og/SxXy
8j8DUdNIVtBrlj+Nq5nfLvrGbIT93yOIlC3J6obh+A/k341O2Lc+jb0XYzkJR2dHieRAmwLs2KDz
5XhsYScHqzubpzv3Yz7xZmhpBlCKr6dxRSOwpDQQ4oNOJIKrJAZWfhW+I+vYE3Bi46Ey2oHz/j3o
950DuxQb1XYSaoC8K0MatXNejtPpmwJERbJYIwNUO8G46h9VrafNmo5q3sdUoP3RPprrPYsQEDKJ
zv6bONFW1GBshY4dPbFqMMHuk+6alsoXrCMlFdsgbVG7I0PQMI4meZDrJ0sGMIlTyNzp4n5134/i
Ie6dgwgOZwtGI4ID2is+N4t/NFWUJoIjirqXJfosSUagXm66Fbt/lVIXZ8z6sha6CnXikAO93juI
/YOgEQtwDNNTyueTjsX3wEbn2I3iCVJfJpoUxe0fuPC34D+8AFhvB5xr15isDTYKuuW6anbSQITK
jU2gJw/N3CNaip0ECfMDTeIQO+5TZxeYGmYTMYyZbt9uqVP5Q2i0krw8NwR1bJx/8G4HE1+ef3cl
l0GKyBzn3MpOukvIV3lC/ZTe+UPLIT5RUnIySWaA1DCpvDB4sXfx9E6AagZvqZoS/JV5uVF11cy7
XFJ/0XTD0qVMnLuop0wyiLo5Sur/OWNccHsQPjDyGj6kNe/0QKLKuNxBcU4q1AsrA6HP/RoNKurV
m6WISq9+/Nk1IKxeG+KevzyMN79KmNs4RSVtWdAS2CV7yJZ2XJ1bHaAfG2dpxbKH90qWA6IsRoGM
EOBVqOozl8/4N5xdVMI54fT4OyDw6HouxFXhJHYqBhlngoM9U01ALdLjdDUtw1FBxPl9hEZHG4tU
tYOBqi/VbiWjSyBWT8zu+hTBK3EBJ1zM3YcX6rFiWYpC8pO6dcJyUbePZWyNX1KsSWiCf5uoAMGY
h464dgHPbXuICvx6RCEy7iTInUx1v5W+fMbyUBGPmzs1/52PmZ/musbeEmtx1YJEHGDuVnE5jktU
SoaCQYPNfa6+iLSZkPgSmshfC+9MGNHBYtOIru85HVRstz8SvGurffFuKu4quxy2laRSVStL9+pB
HNbWIZmtYQATM1gCDrP0SHpLAPFx0zQi0mAotinHfTNaANTwVoGvCeg8MJ/jqTvkZCCkmD6wNjQG
QL9digCe1eBOG+phfrkEgM1ldw5SaZPL2hPiiXUF6GwDyRMfbHuXGGMvUmVmSt2qAUCZDGsJp75o
LzyhAzG4tdZU8uMjyQleXEIeXspvyD3Xmg9A0/QrWmHDms6+iaO/c4y1DP0GmC+SCW/ZxgoZByLU
9Y4XuLNvCYpxRyCBS9/gqH26V/kYGgx2emywBdbr/0bCjQDbBZrtuiCPrB4nrTN0sI6uMRV+ZQS6
FIL25qV2z2iERxUtl1cyf+wVaYCwJTWGM5AnaxE1RvH0o41BdbNLAgMPNhLMfaLRAxe+BEqIrLV8
tADZ/ph2/W5byN5adVOcbdcXaMdUOSRsr6gGU+d7jMo1NoZv4zBLOA25JwESWDJLKLUT+G4aPaTk
VClmu6vF8m9I7y6Je3zNqjVC1oQUrnh0DJrMSNmuZOPljmHYMo6m2QEFUUtBzWnPWizGGUQ+rjUD
KL5R8fq80wKtySODEIHD8elrjKkZP4pBGxAvIkiK8YzYmZcY/LaI36CYRdV7OxPcqzOUSMIk+oou
PJmGEz9fq7QEdOFkgthkXqr121DG0Ech7+HyhkSprHKFBbhPJuuuipZ3mMEHmML4Zq8vkmD7rQFv
7/I2t9aVfBeOHsWlYD9I1Nzh7Pm4k1iDlKdhn8TnJerR9p5LbdoC91xcoLxi8F4WyA7AoAnrM1hJ
O61UkANwiSlZb1ZYv96Gz2IIESjWbWvvBOMy4awUoAFLavLwjqtYgc2gzIyEUX4Zfp7xTAchWhj0
XXVOUmlCWG2ydTms/Yti8OVBc3Uy9kLlIc2X3lUftk4PHvjRM8cFuRsaSc8KjdARdKG2ldkb0mnE
CJ1jO2R5hoLr7Hhdy7wascvr8tsjKE1QA6CJpAAa6df9ySyNyUDifnKyETrI2k5hrZPSWW2aqKtH
BFcLCqjeRj+/vbTcge0N9VkI5yDA2h57sLN4XK6n1PUha0l4KdSqFD/ho+rlew7Vcg3lMXbskN0x
muUjp0YuI75C6wpTQEpCQQ0fRlKezTG0iYKC51NGYSu9oSSP/Hi30hHLMpNng3x38tHQvYTloXAv
FbnRDZqY7CFl7uCfs9aCz4RYr68ax2eyKPVosoLzLsOoqhfAL55nMD3ZxRv2KSeHnMnAgdekQy7J
0DFltPkz6jAisgEAWv7VdLJwinPRiDRX1QbsbOF4SBERO1HIK4Je0e8Xgv/N86gYOv+yClS9HC4j
lj+n6r25a2RKtQC0JAqixaMpazAM5QBboFRtuFl3QaR5/a5H+pyxLAzpycpJcBZuS1bDhusX4SkG
rgotGtFwdxFcpAwcDs5pFJBXT85ifsYDoDPTWY7CCB2ptlYcBS9/zHaSAzsTlGG/FQ+Jh/HXAd74
tmAytUnwtKWQ2mpbIegISttw4/TPcMWftWEljDTb5kL7Hq137qDD5Q2PIKRRq2h12fhhJMQUzDfg
z7WoeIGMV5q5CQrsPjURJK2YqDcuwa8MmOH6wM2ijFkygUtFywqQcnceeGzugvtldXplfQkBRChu
/QTbsmUGFt7ObW9ZjipOkoRfOyCeNTJteWtdF3Xnvx1VjA2U6MhFSq+uvTpw3HKH4Q6tT6FG5j0P
y+vsBlWmITFQ3i52/uSC/nuMvRvVa8ZTpUqjp488MenfB05/fSaojSzSzxYKyqlAFHuYKgvNKDXB
valdWcmY70gelHIIb6+xMsd0Hit42L7rbn+whEQbLhCdpwsPxH/RtrApJEoNW4YOxqcUzn/sqltM
fCdc/bDU2dtXqWe8FVSLg7GiOKzQ/Uk/BrS3y5Zgn9OZvO112qMHixgcWSyzEWIvjXO/46YhoZ3V
Gqh7Qww32oU/TDlj2/pAkwf8vYwn+nCZivmkIngfeiniqZVlFKI6vWXghxrNsNQi/ztFbIK4WHMl
W517e3QuWACn50IdHNzJ4spxTTCfLbK2dcTfTmpIEixWACzI/JF2+uuSPocHTHZRYbmkIt5Rh9/v
AYz6ok7bG0Q9HdZqJAGzwsg161aUEXe4KY5RfrlYX6c8gkIB1CAVDt93cxsd2kM6ICDBV90SwaFl
H4dGz/e9kGhoSSEur96rKCrSU8FhFqdTVzz1j2F8EbaPeqgSSba4JzOJrcwQHhKlqueuhRQIC4EZ
OjrPFKc6KdIVrqZq1g2l/P7dZle8rokcnS0aCAzS+1dAzd/Vu+O2y5KyX/ixKBxU5qjDdvWuPiaP
N/MEYiZh6C5sEwfv6r+kuV7ZIoPCBfEDiuPJ9F81K7MHA8DC2cA6D8C9+gydV9QOHAvXruS6benv
71q5BVuRapDDjLhOjZVKF4k3Ay0mmxhnhFCusqD6WhvL8rl03Cz+KvaeZ037mlvNPscE+1lUTIft
2jUaRP/mNKirZH7/1bN/V54iL7dc800T3uPmzf49KkHjmEwX98WUu5ssn0XXu/IXAnA3DcX+ZEg+
x+chynfyPT7C4l9SRlUGcG3aJvpFnSezyvWDfOKfY6l3bApmW5ZxCptAgxQ1w0NDHE6oIWqFUceF
/Az5rdHeAtBO9bsgKVW7HyPeO1blOWi72jW91Vojs+rKuAlF0v5NcXl037/8JYem1pmYUQNyqBRK
ixfkwJGjR1Ue3jvXgGM3N6W9Hj12VJI898WUmioUKn8ZQqm3MlD/r/gbF58vzh0wljrumNgd4tvH
A54jfAb15XZRcZ3E4MxONKQdxGK8UDjB4rvNsn2Hj3v6dl5VMDKJsEewv9mSQCO/zQpIYEMPj/CB
YvqsA8G/je6RVqys3annyZaLtZDCgzE+5g3lR3hmGpaiESkiywnu9WJ0ygH0XjYOHvWsedW5bJEZ
QlIYTT2b/kZe/79fE/ryj/JMtYHHKYLS8At2nKDlJI2W3d9EZ5stoEPjsto5GdBnGTPs+HytKeGI
piLzU8t1NoodL6YCIPeNCNoMigbexggQiMFGV67rdjI1NkRQiw3gPZQ1mx2Qj2jWLRwHI4P4yCSJ
Agh4wMTKqWNkYckNaS62pDi4hnSLyE7H8DKEUMMlWB0Ot6ikYn16iXJL/QM/rItCVS6ggfc9Updo
JrKmooS/VuochUO0t0qiekm90hDzoIqnpqK5xqNh/BjlPujsAM5lTO98OnXE1znYCrc0f72sYFZ1
xXR28OZP+lxg9jFxPseYg1WK6s7DJEUCYw2XT+i2MWdMvmFYJFlXR4lOSQ8Y4WoZXKxkeAy9R33A
DPYtYGVggc/yUwbaWaffo+4tKpupErQuGjuu+UoxELMW0v/cYieEYNWwzpxM2fhL2XNhvc2ZvLmo
kCqYQl/GiNsEv35ICtAhSL7FGBtbM89R0q6kzpsDq7VPF1HZ0VGBZ+XEuASjS6QkIiNNQCr7uuQ1
4XzX6gTct1q1pT8aUQz9acOFDKvimjGfqWEzXEMvkm7zROE3r6QErqepZ4x2qIRL9zodYC2MhaT2
9gSN/2ZU6W1sDGqgmYXIHovhkgw9a7Zhj/qXD/HPr3h9JkKRjAViF+MHazcdoLnOKl6YEXINJ6Os
IqIGhpx5lD/kDObGjP4yrIhKp/HBYJ+uO4Jt3eFjmTVJDIUAWdDsXbO1eSAyIIO0xL876MUVW4As
VoxjqCZgYDIDawjng9wULdee3LQ9FrW81VeWotacB4n3gK9vUZDAjAJ6SsV9MUffBmKAIH9cVphC
iibNNCjHH/hra7iq3zbh63T7fKwQDUilViou7Y5ZW3Di8Xfldk81LMXEeKAS0APvoSA68e6778n0
cioZcnKC8DvLWot80qgmkWPYftxLB+Ms1HkvFmWzXmcSZ9zzq8bDQrPymjq+buTZkqq9+iC2/VLP
RBAmjAwfVzQYq0KM/Qlx7LhNKVyBHe6T1pC8sTTZqX9bPtShBrBecvSO/uFfLpivIZjmIqLgeomT
NGmHifK6BaDp0iSDezyAAO1qSdzyNNkLR29YCos2wcqCru106MSg3OjuJmiN+G5sLBwKqnLRK4qc
g/AGWP0o3IebMWGZ8+KzfIbhqmr1v5NtZR4lPNl12BkJWX4eE2R1JueBehRagcSSDOe8oM13rfYG
olCUvtrzNuYzgPkycpGb4Wvh6RJ9A50MuYvnxEerxfSLpeRCBpVdoU1NWui9LfhZmoU0WwToeHDQ
i8uBoe6f9fCL8GCM7JbgD1tQIAm5TUVoTpA7JOJl0FlttUrvUODwgZoxnWTnlByLplX4hwuE0DlE
QXzD9gArAGg/kg+V3zdh1kKwqdUYq38qxsjQoWn7b/a95pbn7SJaZKvt1oA+oyf4S+6ew1CAajps
Ujl0JgEohmtQDxOGH6TGl/BXhMrlrET8FrhZueIa1q0QaziBKR5DncBuSGwuRjfl9HpGbNkcwbDO
tTa+U1n+KXtyBgOoTUSy8EmdyG+mzykQk54MXaGQflhotsjANIzW3yb6zHEoNFA+4QklAxNE5YHd
bhGSXB2FD/LMS2DRsbd1aBIwvIiQVd1IUl7OLfby1JGreFILaZDGbvJQE14+Z4GsvSCPcdqXo1Qe
FxIbp3JNkzTG0njrgGh+LGFwX35dNvXJjr63FLDo+LQby80QqPPUGKU0/8XnCFTNk3pwN2sMIKiX
06i/D9cUu50ZlTcQcbsssg2xBHCdMJF4q/4qD7SBeeqgGhrLt50z8IiEaXoI2rsa3neokU4MoHmw
e5cvvobw0s/M+jelMJd8ZN0mFeuPTsNqZwMMIY9n7Lr3+dq625rLHDqvKuqh0ZaYa7cUR7n0boNm
pPkjBqjlwxCjWhNFrMXfUMLKo2wWBDDb75glfJ6d/LsNUG4vHUrrRD6fc7wW7JpE1q6SOc5RsHMy
dgFwafwnerKBRvrBezzPnwnHhBRv4xQ68cAZYh1CAPV0ZRUNUe96QJBJCcy8a7unu6oFjyEq2jjH
M8HLGmW2dYIlQb0luw6W9yqDjDQyS4gIQhc6theHiJ2G1gA/cKHAB9FATdmbMJJn8/PukQNThrDo
t3eSaJF643XdAf8WG2e6XmfzcflnnM6XhZG7tmAqWxYhEPhihKiYiGOMJAAQks+IMA94N1xhcgv/
u9C1aX+xnXoEfDFipOd5UFgm8iPCaVYkeQ65Gz1YIhwUFLVY0q+c/oT5QfmjGev2008eGQxhMKx+
26VDIDokMCRIo1qRKm9K/zXQpufhgt9ERbgNh5757EWNDpU9iz67iR0ntfb0PuSBoofTFFa4Sn3F
by5wrqI4x6bt9irxvICazrphs76Otie9Q24nAWbLg4/wn7LDHZqeWLdTX12gVJYhvOGYguUqKvnM
SXaR9TqSZTCndPRBC36J9hByF05oRQuYSmTQ4sZvfXdOPv8/9Zj/fAC7rQhXz46bi8abwt8whk5J
9MOAkWjlj8ArtpaliM8snNw4W0QbjB5mR4HlXM2Bo25ewbHeAdzKYg4ifReu3T9YsBgxbcTHMfTq
H0a5elB5InVVkPEZeBWvsbWsNkL/BgDtfSpr9jNQ4dMcXmRMnSP6EjXMuVyjDmh74GJJSX3vR8Sl
SEbpStaF3PuUeqJRzXr8xLvVTo4CNkJfRH3d9R62Y58Fi2p0wuXkV6crTQPdt+uslPWetnNxAlPE
5XGzYiY6G0CKiU5eYjEzDMLHbXz9v7ntDpsF7oulnbBg78PnC4fp2GTwG3Zwjbvg3CP/p3q8WzJQ
Ncu4g0y3IDSk7dJyIb1uTri/4BBtTuxTXxnj8yAIvWvRRsRMITfO14AdCry5dMREVNLjtvAagjgO
BYv6FKMDV/ZULqcnwYL3AkxX3gEqZBea31VlpFT8iCZV8P7gup7hCOVzVJcEP8jEZrzduhK3K+4Q
NktcXxOcgpUm3ylIeYi+nwsTuOCKEpBhLdiCBKs+EPq7Z9ion1mNDoYEoWqLrPsgQ4hA6+EzUjgA
06FHzapUBinmgYuOWXyEmWMYqDTET8zACV5jUGUJZSX/1YTclWNqh8AW05rXwrZ3PttIuNaYOaVt
wF9qPinniQyeC84ni1bwpFOD32fFf/5VLIcOP6b8AmaupMmuSMCJRM1IxoGjkSll5SHb8udtSrKj
Z7I5Po+db9VX52bijiyukizff6z+QWgq22jrMYEWMecAdLRjw8vbTR7GJcmCQhsntlCri2kSmAnN
AbEL7ysVBEwEI0KqVa6pZrlvmkSZWRLnSXWpPpENQt84tQMKoo1vYGjUZyOSQmpTY5KjUVNp+/xz
MqbZydGB1dwqo0qJatsR3GOefK2w3lJmbz9PQ7eUeKoK4TERlrECB4gdQK0uLKX3KryqCbVxyU0C
9lyGLv+r/gemvfg0amVd4xtCr1QHpkhfXr/iQE113wzRZyQYGJ5501S5di8vLsaM/R55yzyeIn1I
ywuHzUcIu/WH7yZFdMWWKMLQXwZ8cbXU0d5NR/a/tXbkMPuV3LyAL+ILTR/q3kZ74R8ULaZ9pDAP
/G2cLHxxQWH09/Wl9hYDqXCHFf8B5ESN6PK/dmYh79JEa1Y2yAF8ddskjVPZ6NnY1P83UYVwZozj
3vmLipaQwuYiwNAdbvFPxoUyxUSWOdCdSiwWcbbH3FktZkD/cc0mrnhpJ/TgLDI8PkAnoB2dU8GT
ymOcbWOfSl2fFlKZgjWXKm7igGpNEDlygtV5Vkim2JAL1Fx3eGLtsgh9DnYQQox3kMLXgAZmkqUz
2czkZKfVCvJzcqyE+qJ5WzRvcrbF6IJP5ajL1AAHECmsvj0fHKp8iU6ihPDsx5jAmPRtCWd3bP85
U6GO053C4EiyP2cnGtudIAAerR9kKlZPw1YGpne19p3+p4VlkHM7gwme7V6ikHwQg2/bPA9L4+2m
veROQya3ebMS3h0SOD37hgGT5DvH/xXpz7wvePQSFigu1tBANr8lO/2FPInHVaqIhJjF0HYBFVBw
dIxTzeaLaeuynhDSTHZU2Gfi5yqV+35Le3bhWUAIgbEmnui3hJDMeTLl9sfEooKziZoli+M3NwPy
EHoW/TuNQ42oW7HYE/32JNNtZW5CbpWET9XCfa0+OX3udtZgkashI3r2BPviEN2j/jRLa/6aKnEw
REEELOysIC7zPEC+bOm0FWKC41OxYhUFsqibrnEhD8w6+zAJoy6Ulfl5ETRs1l62y2qhRyOGLMZi
o1kBMwfQFwhL25MmZAaojXa3Wd5hwgF5dY4buIGA5sW4QhxfQrQzHQSRo+oWlvUXKPq5kbNUCqRR
QAirFC1ntbGx5+mcH16HJN2lSFL+PfpKBodhHsyMAEHQJOIRo/uSmKKA+PZbZ/+nAeK2ikoEVaFa
ovvHKBHLzUoO1FfPMKdiQh3nMJPt8ZIfp707OgjkcQy5Vuf6vu+d0cD/yGV2nfMSzI8QruYajgx/
OJMw+7Cy5S3qHt/jD6ZvnHcs/wkVLt3eAuBdZvuwKmXfpVcFxF3iYq0zS92yH42gTa+PRTuBQrSp
BE/oUI3NgiEuWhagAWyY1PSM6pEV0pqOG23PGPB0/EONklqzZsYNb+SE6iDvfDLcRLsQ5EzNnHU8
DQFB55D09EZn7pOIXYLAQjPh0jTtj9npFLJ8K0D8I+zcGZehixu+9L7VWiyiob2Fuj+JTqMZw90r
ZG4wEGLc/CuVcoc4OeJgd3MDPPWcfeA7AVSnkb9UHfBP4m5sglngh2BhZ6fCUFXZZ2d8Z4WRwkfv
SyN9axfnM7V5F3BnCT70DYk/7oThF8ad/iw+5MM5OHlN3S1xQr1Dm0KRtZDkUsTEN+l8rS1SwipI
0u9gMvBkykUNMuATMvV78J7BVYh5qC8hz/ln83mNH57JTZBzM/xjVYhxhPYrlcF4Dtvb5FbZ3Cv9
+tlIKiVZmNnBHPQVB8Mbgwq+Ox4atULSbus7cl8FBifxBbyU+mXh98txKu2+Ld8I1G+aZ4VLB5oi
9H/TtTXmq4LXtCnK3YJarbMq6bAh1m3q52CxYDstyjwgsS3YGcYIfQ/yyaKz/4NgVoMlZWuUrciY
5/1HM5Ep2/mg6aa3typArXi4S3QISWbDZ9Za0yjZGpKW9M3Ae7W4mjSPbEKpZnOseco265x4XViB
b0Y+ZvgZ6RhHqO8WN9QmAua11DQcMLPSnLh7UxkKBRARBMCjGxxzaOyM/uqHsLc/0eMYTKxdu9Io
5QKFcy0lskgj1fOGqzKcIn9LBG+GCPP6AxyNX38voYI3gNpiG0fQQyUsqn/Y2ISsN96ZAm1yYXt7
5HKA5Lv+ni+KN3/GwWITReJuiVUOt04dRR4OCuaUvY0RG0OgRvGR0BepLaR1ctn+oLN0GfDPBNHR
hGiVFry2XzaGMdz4i8NyrFf8UFqWXrUAWd+sV5uz0JzxzrFArCZnZhkdiGk2saHKb4iXD0xtM3Fi
4bPVM0J3jHVXcKhZZO7ATT9gS8OeUyzDMDFXXS24omBIwx2DOw5TEQvrx0LjPPL3ddLWFltXwBSx
k/WuZb8EmfKNS1LolCFomlbsctsn/FdBQu04KDCPrCjW3Mn+AZg8YGd3EHkWcZGERX3x3cX9jx/U
YuJeQLdpWz+TCZinJoZKIqrLW5k7NKVkUXV0fCJIBUdnuL3tFZh0XBB5r5i1viZHQW3mxr5UnEn2
KeHhFjD/kQ2N90PExZ1JLuskKofPQ6L1c1a9PHO3xZluEynD7fOcssBUewqH00/YUbLIJ0uedP5P
2RdxK82Fv05j/1xSwPzojCCRwkdlmXXhbLtaDAmz5AZeplJ/XeludkjaKnqCvWSUYp4Ul4L8HgUm
l74SsyHmJLCs52vCxN9kKWL4xR3l3Zxbbqr4EFED5rrgx1Am5jopzWKWJF1h9GbJ1SPh9g0rY1MF
uCOlCRLcV7EO0mi6vMsyYE+JE764WM2hBV9wgFqaB8RbYdaUynixVNPah5oT64usNbgSqe6BkI95
M2dGnD+Q9OE1BffigtBkSSbvwgaLs8qH0yXVJdfrlPtXvQnRyeeOq5doXpS+LAeRLafqfBlaDkrV
Q9YKP87kqVWKbd5okE43zpD7LCuOv+oMnlvaEgMPIJCabjBL5BNIWxdiGix5QcPJ+8eVADpeY+S7
1KY3Mhr9i0h44Ghj9DdrbBU0vkINo2wpj/ODmH1w0shPUD0CRfMcWuqQrh7BsP1cGngHwvs30/FR
NkBwQccwMgPKAEZTjPFTHTSKkT/aT4nU5vJCZF0rK2/1r65eGwgTIg9NEaqMbqB0pUVUgef+K9wk
g2qDGCu4W4vrzIcWzBSUe5Df0wpiqIN5ZLwb4TnYmZ8MJrENX0fy5msfAUwD+af9YLLHAenQcHDG
2a9A6lFvIgm6/wwe93D/idbMYWTAufEdiamtMEMczjHlV0mqJV0XMDIvUU0x+8ICxfEfU6kfpVNh
GCWdlBtudMBeWbQ+xy1HZ+vpwQnIBoTAfYEcH9ZUtUJOlqWJ/7a/IHHzBZt2r8e/N3tNJdYO+0+D
N4u+UU0yId8pdaFZst1WeCi4uzQwxm/auW43rcpWYCtPwnYD2U3EDL6bwe2/y0ogEWYDEf4T/bDS
sW64j1nbtHXQ5SQrCkJL42tWkjPf/R17VuDFzqos9Q9Ycemaa2vofOLXmAKFpKEQrtIfjxQrgDP2
3qBRSHsPLL8x0+aa31Ucldo2sRFyxFBrCWeFycr3YKTFmpEYD8FMD2Dtgc/MWKPAGtbSqTw+ybad
hUu9LXQ/LwT3lPz3d5OUya12WKaqmUWozdlEQ7GtOZ3//X/RaQE2W1f7fYqP4FLjP8ACm+x+h+S/
qss9UDPppeSEwiUnxlanm03elpAeaXj1T4FLMKGNMou939JvK+jl8cju+suKXBFOODfcO3AUSm5L
qt1af4lZNPd5HSB3rZ3KVs+ZO/Pv//TB1ErJ+UF3btF7TPyiQAleerQ0bITQRt4XdXIpC4tDXy48
cU3fy13CtRI21mS/nOgtyxVVlG4TP0CiDmFlFJ+bdYXwTO/iRZ3984ovFX0QoPt9vWRiT5CibmQp
mwJ1ta8oGKIx0aaLrOrnXgRVMpWtMVlyAxTblZoApSt3iOeDMRb+kQOvDM3Fm5x3yIBJQqpkjzVI
fwWWtSxQpxhENcR9qPjqaoosKGFBqOy46ONpWhsVp149seTBgL33ZImFRSEjyuxpklsOYJvxIgkJ
fsBtq1gG0gbAq/JjeYZqzWA+zyXlgmVQgoFKUAvmLG3otVb6V6exuk5t8edrc0SzCGdutemEwl7f
w7GXXIM3Wl6F7iPfHnESAcfWC1Kzxg4NyQYBeBeVkWyGJVR0RnjJr/wykt7/axRJiY65Q14MAA0O
+zcO5TZ6Qw9nDm9Le13M3BTXKtQ3jqD+EgmTBCI2m3twyhq0znhRqr6HpW1OKKqNfoZUDp/RXTy2
0uXIObNNbOY0V8iYihQwbtR7CCe6BKZSyRMNP8X1UNLaUCLsHQYWHWzHZSV1hhsOAZYjGJc1I3ty
8qPFX6cMl5J3qTJ7EsmpAYfPq4JcRp398EpvA4JysiEzzM4jOmqO13+OOeNzE58wWQxwi6sLwDPM
bEDoGPdCWKWdnoD8T2Xu7FbDn0NCrQTbvnDT48Y3YISi7pcLCg5mKi905s7fqV0GQnfcQxrIyF4j
IAoGf3+DcFaBDDN9cEpZRSVZ9d2/UZ4nXFVnmKZt3Z1eIcBuevwz6gBB+jAsv/xTXR3/LZBGJfsB
YPqtsMmMUP0yNoAttkZL5rXwlGd3RQF2MAGYs5e3pL8jyowF+a5BOQbVcadWMr2hZIMU1m2RQYqh
AF7EssWFjHTb+L/2MVw/Fd0jIK3TW2+1G6XLZc3r9fcCz0vW0xj3ew6dMZw2+CwlF/z32k2UrWOn
r9G6AZVR2z4vxM0gR5OMh3RinMAb003WQSq3Qyq8ibniH/z2PopAOHNimW+3K5N0jhKZcu3DXW1z
8r3zsZs2QosdqJUflqCLg26bvJvQif1RXpts3JlIS8EUPlATBQWo/hjrxXhPyPRLXCHVebWI2asL
asUQozc75LR8T8YUd72lGMwXoJfRcku2fG2ks8NLcVWrvUewYa774XYtni8x1sjw/uvgu9dNERgg
15t/CkB60NdYpBKGkmEdCpp6B8cRx2X3CCuoQD5Sj9QbOzNm29MQ9NCCiweJShrTcEUax9q2KTDn
DZKm3jlJqZ1Tq4eM5ND28GNxp+7zjmt7nK9ysghN7NSzjaEoeAPWSQvLBJvo5N23B+hZWPdtRcgg
2vBLLfvafUoqfQl+Ov1+zR1V7vNfiUb+foE+WDrx4kCZ809czy9R+cAe/F0LmadFSzlSD697Kffw
L31LZ9nb8yie+QO8hC/LgDGNpNz1OjO9ot8CXDNY8Yi3VJQyz+Umdz5of9jxu+yS3+kk4tdhs8FD
TKD8nvE1k8Q/hTqKx+BaQbkDotPYRLZpouhbvGgjTLWRCdII8pekK3IGspf9XmUINeD44LAPjsLb
/YdWxVYBlrJOinqEMm4oykoavmrBfBcbJ+ow2ODzgtLcvbdcpVY8CTDN3dt8EbI4HlxFUlFU4dD/
AixjgrOwiduuympOu1VVdfAN8HmbBC/1Nc/Ts8MvFDGQF/peMdd5q1kl90oMMFE/dLsIbR23a6ab
zF12OqlJC2waS1DCzZiThMeWFBtaGEESAKUI6GXWDIyCgbGRqNeT9dGj1e2Ldxc2c7qUPEFspTHw
c2JouVtrZvtm/au7DoaG1Q46nJHp1J7pkmD1+s0P+UqjnvyEILVVLea5K0mnRAAo9CDQMASDvxuV
/4DWtUd1T2UIMG+gnu5ThKCGjP8B7Ap+rWyoBWI6ZhSCwF14gHJ+P3vYTGKz5uHpV77AQSawwI1F
X8ji6pKPzWkaNB73KFSk+pQNjRFni7L7vCXJeHpesFuZBPg4Cigtxu+6/PTXRJNsWoZGRUQGb+zc
gp9nUmBeOrnBwHpv5L4WtCYj6lekrGGNU+MMb16IVvIeGfrYSSK4B7FzramTaZNkxZR5mXB/4bOR
9L/mjxV+FxBYqFBlS4bBpy7WJjIhgi/japujmkQssehNJDZ379zqXZtjAP3kob9+n7aQ5vnvfzjD
qZWQts+EUIFM3w9AmSedtOZ+RRPCMjgXcmGVvBRHP204GYlHGwJafzrFIO7GxyGPFe3AsAOx37Nz
NXTrAAwjkk8GNSt6flqcEJlzKF0BCIB/Sl5fKXMm05GdRVvOA8Df/v40W815LYG6tVrJ52NHrR2m
OUVFhMA/Bd9gwOxaRqY6OWe1DXkP4eY/fuJzyJAogB7NJl16tlDTl8GthtrGuaSXapK/SeaDBPHW
ay27NYZvS/YCJDmC0AfXBWFsw3GpTnozexJfIbk20KYXBaAL34YlzmoGEVbw1NFrCf3rxwQ6eYE2
B+7aC0NG5ZwNLqq9KpLpOd0ehdda1qazAoaRjysxHBdaSpy7hPIdURgcMNQ/m4P1Erz7MdiPo1Ml
GlwS6TgF7EX5ykZ8Hb+x9wT7lOmLUCiqHwrwgS8D6dqpn8WQUpSGGKdHwR7FrbwaXYTGJRXQl0+Y
mqAdPnGaLRQejTdNoy6wS2CUPc+B7KW7RDSoI34EqWl+fVmxuIDIe2vikJGyk+SEVr60PxwVhAm3
B1xUA3kpedoF3OkWg3AB5g6K4YbUOqO/Tmv9tREr2tO+T7slBM32ZNTw4T7ijr4WJyS9uK4YeIXo
1Fe7Agqto0f5AFZZMRScmrns4fvz/uXh9+OQCxJDPsc5HQLW+CgR9MIrTchWDExSs8QtPpVBlovH
kwteA+TrJu0r7DUxRgq1AMLi2O5OIQwGCGsomSIoZyk+hAoCyFzvpxzNS0pTK/iUOeFSLOiPD4AG
S373cqBl5bY82pe5RveCw/XnS5JP2pGI1WZGAjI9mDtS7xxQw8BmWdEN9qBoFUu5MSNe3LeG60zl
DhQNCQMVcbmQX6VqbkLNlhtM863t67MP2fUMwgDlPTFDob4tllXVU6vAVoixSO/4xnaBNK71jCMM
Cc9DvCQd7IjoKKg3MEjAn5d1UcZDobIDndLMsNBNx+u+ULnTQ3YaR9jhzdSWzhnB0eAs8UxZNEpr
gbSTfhANkoe42DZnc5unoy4ayO/sGeeXDFrVp24g2YPiO2Fas88r5ttu2IwdV2wZiRdGxObno+vP
2b0Mc5W5GPbR/WX8PgH+WaqNgewVhALSh9uuRiZ8XO/1XXYlG2BTbKUCy9CZPAZc4yqARHLoeg5g
bbKdS9pgCbdtHWqOmICzkNXYOyP/1yLsX9iCLqAQ60Yd/CAgIE2sgQOdBsJkm1fH68kSmqJs34Tz
3icivJ07MDzBEY25fWMUMXyt57BJxAHWc2x+wagp5eFS6fEIQoaMRgtWFyg9V//3mdmBMKrEIzYe
B1k5/qxpm2XThIggv5lp+hN0FOFhxbeB0MP3z25dW0C/8okeXR5vM/N7B2RAQVDVOHSgKOM4olBO
YQCHa/cESLRF7Ao7ZyuipOyt0gtW9swbDzf6ZLoN0AI9PfyAslLVfCkV03kWNetjKTRCyd5eduMd
AJWI6ZkIGVDHOy5FJyDq1Sh68L5RJ0VF+Ei1eVd8S3HYFo7GAapJ7g5pKhj/uI6NB3RMzP2BAlwx
hgK5JjfdbwYaL5a0K3c0za5NoCHxZ0gVxPv6oBIqG8I1yz9xYlOb9gPAYn7WHsvF/tkDqKxkjBFW
lixtZuamE0j3ftrnpal7fKCtTyHqhjMbV6Z/IJ967l2/EAoerBadq3rLOnsLWZoOpn57Csn0pgVb
sba5I3s80rO1epTKs76h2W8rpjHkf9M2k4phV27nhZqUqphNPXbQAqok422hB4Q9ReFgXc0PHSmT
FyBtBdYWEid5e3/DGEHyuVmOv/AHjWo8HXwBu/Cg3HezNdwDuz/XSDYmKaNVdK+A3nPuGJULDl5U
A3oFMq1aFE/B2WDr5yVt/xz9Coe0Opu250XTcWI0albgRBprFGPSipj8QqSSQQ5Tns/ZUsDnC5gO
mhq1KbODtK/kPqkIbe7me4LqYJe/oF4yZc2CU+/OuiNo5PxptQ3h/0B/B/0Ayf/PTIRFcvU0b9jv
EH2ECAQxXyvjcB+4RIu1Uh3W4q7UxIUoz4s4FSekLhlVBlYpXowUns18jHc2qSkEZSsNY3XdjUZ2
/kjmk6rbI4mJ2L4Eewkk8xyIInce2WRkq66Z45TV5Nn1PwXEKElMCs6BVQynKmusXeCMVhKeQoRd
sB0qinOFz/s/Ctc+wyYwc7DiJHG4xltPOiBw6XQZniXOuVxsuOU+Ja5qSaHVYUz9hMdhR7sE25YP
tgeEBHg6FsR+hf8+2lQFC4MCbFecrpkDyw2EG5MR0nxOyqgrDM58HfcuReIiddJzBglOX4Qg5Th5
Vf8wLqoaBofeNe8Mkh4qggEwOVNlhbieNR/Y7oPd3Yk2yQPxYIIz/f4netKypFFp6WEn5UMl/k+j
7BCJwCi4oSYVWcrOhdXZosuzCgzpAF4bP0DLefOeCvZ5TqXlBdifoEY9jN7vJfH6egNEjUGs4khf
S5lU48HgLwhbltHZpILgHg9nOroFpGZAtUqklvEI4rmxaf4OIxiK7foeL0gxlR4t6NKBWxmKWqT7
np7O2rgBfUakKq+nCRai+l3wJ8iIhwYiOuBEGlkdzWNhUiGW0iWSQLYKlde+85cwifBtq8wj0zZp
tCw9efwLZiH9wv3yMTQtTitCpgUFdyEVRqwWVI5ykhy6ey9s+Grs+yWCrrQmYNp35lJgv/1I8X3g
aa+gRTNrR5Is0FDikj94iKKjwgicC79dwG8EsTF7S8Svyi9Ku5goyBjjdu4ta1u+fi4As5URsew+
fZJdFfBz0LdwIW69GaEGvFfXTWdwenU+aQoSClKGwnRkN2pdpLrV6R5NAMODHB8O6X94Ih26sbdC
tXhT5UXxaCQaGciytPTc0dkIJlhV7HfDfAu2JUIIYhsAjqPDvKRm0Smzd9E9cttqrNEABkDQNM2T
StMtSkrjCULuqGDfrY9mne2GySh7pXLMQ0oVSl4/61vFB0gmnhNQ28aYFzjyUnGVB3x4mny3TtdT
kYgKIsW9IJ/nO8LZ1SXwi/zVMdblH0lCWy8TtNtYhx/zjLct9fLXB3mubdXrRtPDd5ChqMaW20oQ
PBbbZRQ4jN+qjRUkA6rmTfZKV5VFauuxndgtokeCxlveGZ5KTIbxBFER78btksFbWBOO7DAm5QxE
4QGYrzA5QM2+NxG/LjEWiLvIxcMXxKfgwMqS9ad5A9A/LwIzog5y4Evb1DnS9wI/AWZvEjLR3K7O
AGrtk79I+bYctU/OG2kK9WZ9PeJTBYWiKLiGpJfUDij/P6UgunBZmsuWS0XWj5qJKdNsq1y+JSTY
ohQkbbs4un9JsVr7S2P2z40lC4ONYPvr7LcJIFlnjy4272ppa6uP4+zJjQdiLQmZErvvCeDCiWaq
nODTb4MO05gJIXHbW1hHwayYaJEVPqiNLDXSmTFFWSg3djVrEQ4T8QMnDb3KBmu9zYgQkQoKAk7/
nbf7xb0TottKm435KZkgtMpx5jZeb2pltxQKJKXZvua9USCSGF8b7n8ZTLuWsxcAeBYr37v2EZeI
rej9pCN5GQwOY3GAyo4vjyB8xELTuFz08GZdiD5/ZdB3DoRcqmATayJSeYTyf88AVNYxIjxacbb6
UOxDXnrlHME9KKrMI0lLOTd1WWRZuuoJYJ9a9bNNkiMjtT+vYFWDX8+iSQMqXzWFBzmyo8hBvQey
JwwP93AatUv6g0My430g84enkCLd1SbheVo12lA+lahbv19/9yw2NX2LDufkynLYTeYSG3p6/Tf4
u2KzF7M3iK+SCZI96K3xb/kvtrJkb5j/Qmj4/QY3ulbhCTKuT5AIMMWvMU2D1yA0i3JYeqoEir6g
JhS2DX+N5S2Z/7uJErYBcG/I5UqcFTE5knHDoh7lKlwVIyVD6TAlxlMBC0JcpH/5QISLhHTiZaaw
YSYLFoKCZhSw2C+qdbhyPkSaBv+TTfwvZGccDLTVQmrbsXsfSQVla1aRBhLhKBZOr450pIXZ+s6J
zO7Ck4f/iR2ahiouwiG9q8TK22jdlaqBfRkYu6J6ltzCqg77pVEF9gCmrgF00sr7CMla8Ux1Yj/c
bp5Id+sPwhBeLMl/ZAoz3SPsosuzKwz0Mm4Xs+WYIH5Le5IBLz1wJ2wUL096TF22KDLpuWsd3FlK
Kb3oRmooptJ1OaNEB9vU7C9D0DHhY97Tm9r5msuzuVu9/4VCurm+d6BXad1IsPDFdD3dOUiaERz9
1g9cdnhBHCLXxpSDGoBavQY8PxGcXgkZ3FPq5cmstArsUGWU8aaNgH4yjQvawrxlNLvZtniFOXVa
NlPry7GKIyaWa3GelAhDvhVYKaNSSM7tYTEu3o6VeX/MyFVUZgUh6/gMDFb8hZuwtmOeyqw6amqC
1N2+HLuwVXE/U1rZwKAD0cTDfSgoUwSgLw/rgotkj2XDe0DaWxuPxPo6KFcOSj6cj6Y3kl13f9VU
PkZwJ8uU80MWxQ3jMXUrOwpA2ohikd3IiooWQK/qnLX6BVv+OblKXUdOf+mqvzO2GnXFw/dHnnXb
OkPJf/QC15yOXL4Wp6qVFns4tnzWIDj6xtwcNOW6LcTOnTdFO7xdS6rRFVB1ICwmjaAbB78fULkE
YvS86aAGlbxRnTRNrrE34Lx0B5qO5Byfw9xYGUeRrnkYLwotWrCt1LqpP5+Hn5F1gcBVaGrAe22d
Bo4g6DG65KZy6nufk2SQlPUit9sQs/z8bXMEwkX7c2jShvSXOHBEnSn4hgbRHTlqeKOtfjH4ZyBd
fEW8EoYbVMV5O7c6ssMHPIHdfVfkm9qlzpXhDQlvFiEfTGsa3m54JdS7vVsXDLF5IZDfUOQTtqZx
5nPX86KTH6AKCrsVDwZOKIwLHmcGBtkLb5O1/pgUw1wa/PVeh8reDjYy+poBMc8PhuDYScmAnA5/
qCd1ZGkjEEGKWxfx6MEFDk7fJouA9JmzDbD/hdit3u193FM5Z0AA2G3Au0dLxMSNESyxzB7Hmhm8
v1LK+mUxqJABg7TgaKgCgx2ahBjQb/VV83pFlFbi3+wvWrO+QXtZhRYREZg1Zg7Nn4xcFCo+roe/
wdmMlL+kEQnQxPGn5sH/4G3f8haCA18nCS8WEtDpCOLLRQ0YXlwHlcpfd3IIb0WD9Yf9bXxlEb2Y
w0k21OnSgZ0FjCZnmppFNj45LfA/kmkqzafxExIkAJ0MOPcIE5pG4Hd1fW1Psgnme2a2JKI3IoDM
H+v/DWrEKduMmOmuKs3BssHBB6T2U3uqpvLaP/iVSRhTTrI0Fr+Xc3m7WR4hQy6D4WMwP90JJe6a
qj6oJg/kpjXzQ2q2xhmOaY+LkxOZ0PbDfc1ZAvwfV1nt9tumHr4AihOI7wSC2lXG779qxQUeBb18
yonUA8AhtH7ivEXbyPvRwrtfbmhU5+hb5Lm4kaprLJxcNgJv6cd5+B958mkNf7D+YHLyD35bS5y/
c89vKipqVoEh1KvMa1UzKtiyeNJBmUP+DLHBE3fXukL4Gd5hcEgu95im6DHbqpwrT7u7d/pemJlZ
PEpyM5NeFVYCf3w2B5VWeMUpwDt+QKteDvqzC5rovpZsFHyBiIGJcqL9NWpJlTwPMwiKVJbQ0Ctu
KhQ0YTQJz4LGdJNfAqhdAryt9Glii/bSGor4Sd6Dn8z64TCk+l5B44AKuZnWw7xg/9Jd7iziwGLm
QXit7BD1SP047LqS6jgofNp0LfMJzPXKAVivo6X+9CKB+CNElGxSQLzqco25Ou0BN1goT+P72Xy9
pnerHvWYy2LQibROWwjibOH3bNaYHobOk3UwU20dqD6NETGlPiaxyNR8yDlYT7jPTW3yGu4+bUhJ
M4hUtDD30n5prYCGi85OfslARmVJjUXbBQP5XZBX6fdLLnIb1zIElPUvtFRLNstG/1AO1mp9UJeE
ugbbI4doE7lkPpuci7Jch5aGdaBJ85c8VAcQSWzWBRHFpbWNG86oH/7qpV1om+Im+q2mwbMD0JZZ
/77sDAr9BXtWAyGbnEIVByZaDeslu5DEmVKRxpuGHGbHcfm9fb0WnjtoUJ4uujxQ0iRI7bW9dcx+
XArk8x8awzjLqUlV3eyCs+UjqA8kwu0QIkNiYADcQDLD5/SWGnwM54ayDVJEn2YjCxMnSYakBoNu
Y+hnIZPcjQRKo+fYa7+eQ1RPxqj947C38Fu+KZpdhj37RSY8SUriLyAs/MDoBElfwif8DbT9DGhG
hetiV6KSqiV666xd3bpQC0IDRXB6eRYPmVWdSxs9xk++ALSab6dOyjMW+X5XId4S36KNhqTTpu60
btUMTitVdGwgW6SJfWUkf6UoGAGCH0B5gk+1uaNN9c0FuB87z7t54LuO8pBktn50esyKZ+BClrk4
ZoM024Lp7WRvH7UuPLWZ++LLvi4fZZz25gz9oLKtZDRBMJgQowx/AUZkw1BD8rE4DzFydKtHBux2
7A6jtlqeISpLFRP6gvd3wFi5EmrTCur48chh715+2yU/XM1XNhev0LAGLF/BM61WSpMVfGcxRil3
DZ//U5IKPb2vkO4cnYQ7mAh+BYfols5zc0QEA9CXXPlbeXWOJyHmjTfFZqLCd3AfGgdAXylkHns4
6juxFChGFxm5GU3zkgKWKEPAk4y8tsG3uXNa79HEcOUweU83hFbZzQ6uJ1XPLFPaMQytTA+bxgXi
ppOa3yc+YN4r+l3cZ98Ue9M9LWs31Ry/NAwhD0hclwUEo9P+4Vr0Sb0Joh+BS7vc+a2DjZdICSxH
j3VPneOIHnj3scffiAld32DEFityxfEcr3c8q/yUD0betTwrrLRkFCGgENdgJVtjz970cWR8C5MR
JOONSDpXOej7Zine4nf6OHwTTT4s6kx0FlA4c/N5pfXgWPXJB447nq1P6ixFVzJa0bY3911zt502
5d6bA2XkOLdnHHpcQ/mDPikRecIoD8m2DtMTP6/AvfldVgVpr4KsNUnpDDeEBY13hpKZt234iozu
QoPg/1t5fdGwThFpl3aQHr/jIoKt3/PkPHi8rUK/ZI539MclzCi+TthaKqYTQAFHX9IAjPacCB6V
wTG2B+KwXnXTuRsLLWdw5UdBSg8ydnyrS+YTnTRA0pU9qIByDQBgM9Y+/3g61eKtokfdNpNvKOVg
aifoqS8kSJo4iav+ceMx0OVHq8qQY7J5rpLSLkj4CR7IwplkbPzex0GUpmbxggm9N6hfSU8p5vWQ
0qyb4H/3HZS899VF/ZDBbie7B/+hoYvy9Un8TQFWRP7FX4Xixz8nDwIh1TMLTPbw6kWXSRHS73ac
2EQEX4gMrfr+sMt4CaHrvBvXIYGbNCCz3KBjme15kGwAFFNkP3yMCUkdkkUAF8hmVb/W6iv7tvQo
EnDEnNxKN6i8kPw6UXE358CLepCjHAT0rDPH85KbT15RV6WuXbTWWqf5BmSlwIbAXFpjh5qgPcFS
7RAQTEoNI9lZohif7iaF0Jh06nm0b4rHQ7aDIxYvEYJi7a48UqTsMxmz75NuhsvkilJxhOPwlBuF
AjyRLYmX7jxlkS32JoOSX4OFqjZ4qlUaOmIgBgY1e0pc0+EDPr4StYkK/8rQR5n9SZaiXVu9IqoA
jkmHHcbjjq71DFEM1Mygh+aeYfQuwN7o1qbXFTJYgQ3nVLWlbZzjz4je3wsB8BzbYIy9PkypGzks
DtB4iy6blyFdcPnkDBchW5hIkYfFhGRhoD+SZLgV4sBzWfLtH+bmI/mTQ7X5C81j6QcOjG9bqiAj
Xgsw2X46DZ2xEkhgfCfvG5g7U1QT/+bo1lpjiuqzIWJGz1vUmkht212sl97aLTiHpdu24TtBCRjm
5AU/zNeDDXUpTe9hUsgs6888eBxKUvYJVxzc7NtR8D/VUeW9X/qcQDsF5yVNznGU57W8Iw93FG37
gCJerMLAw5MOCvcx9/7FdOMaJJcrTQ3ScL2DdoLlzGEPkuaW+zx3yfSCVB1eDiaAsllnSwaUhaOo
PrmXaAecMT9fdQt29FVMHQVFa9zL1MWb/ubCbpgEN/9baw+BgCEGEWX+TNfc0Rfd4vBrlLUKzqL+
d0QeumOU/M6Z3HOrdyrjpxeHFaZu0oKv2FLCJxq8P0COeFBCShrNkXT4DB6phLVhpZyR4Neo/czZ
hNKU8uwKRbI+cBnK0oJYRZ7XS83Fssth8QvCnOsSUr2fVUcazxPwFsDthRuYW4Is49dpAIBTu1jE
PDEX2coX3VgeZlQV3uAuLmWja+ArfuRUplDQtpQ4l480RTshL2kM5s3cBWg1cevI7U5cPVt0AOL8
EPPM9ikc/pxY6nBTxoFFxtbrWaTojtgNnf/8e3VVWX34dNH5Al4qLlAEv7OsrMBHgzMdrpfHz7xG
02KmvGaaFFrJ0bY+cQwt8tK/dhUglQ27Y7BNRWweklzG5m992lODKnFcXubBfc5sphsc+2YbDUZy
FlfBZURuTEnXFMoW3NA8UFU1sx8hewtYkrC9djMqzASWgtNecKeOkgpYnnjO0w5VhrydZlK0Tr6L
Pq86VE6s/IT9PP4+bSF2fJWSK3sIeUSHMpcp/sNDZciFez+rVqWADrTqdo8xUFUEK4V0855LiLd2
mscK58Y9tFKWtjmK1GDPIdrrjkZXgTIQsY6JLh2Y0fcCozQXQUNIKl6JrVD8gVgnJKvOPCgK3E91
7o2tnMN69RdBYuQf8l2SRmc5+ux7AQFXlfra7qwZrVjzDLS2FpiKMCsbthE2Tin0EbjIXy4U71Ka
Y4tgMnI8JE6yp869o+5nrHcHVLFcToBWRRGjIwk6NPuBvH/WkJQikBisL6Qs8fxIZ27UbOekAaAc
WxmhFbMqFQokQ9YPsQe+j5yhlkAD/LiZYDfiNB6cjz/0ka+64x7pdtM5UjDFHTEzXsvSrY6H0IXO
lS4/JysEc6lo7IPQMhuGkhB6A2ZwIgQuE5CYYdX8g2kTzCu7FMLJmGhRlxX4mDQoAYV5cpgcwj++
pJ/O9l7XcNQLr/7DILSAaxTauH815a3ayFoQCb4+oCEUjtNrPREakuNxucZyVDNwzu7mPZVTdUjz
pJwkrue8AxUmYGiFhz4Cf0iLXbNpeLMfo23K27nQ//OvD0BHQeC9ukl003F41fWWZ3e2xEXM0mrj
ZhBD2XMwiIX/WWQ3ntwgpJJK2M4rAHtqvQtbbq3aTdR0yRx1vB3GunpmeFcBx64p5d/rA4EQlY3z
5sGpdt7lMHBsHuuRV4NAgQAPgYGlcZRGXNFhjt64O9m+OU4kN6Ja5OMjkSGt+nr344dnOgrZ5/ai
pPRt5bVlzrHCcLOzh0D8Ly2KbojlV5kPyERYJjGZ0RMokkVEo+WBvkd4A55Rcg/CJXXt3y1ZM2Lh
/qtdYisLM5VfttrOhk6k52tPijqocJjdSfevhwwFvtNazD452y/qZIgC8Ig9yLuFROKVFFCkLeUJ
WnbDuIHf+0G78Od6DXwOSMoj4q7PGb8Sdp1qpIL8qUwadbUxhP0Abd+F0rPIa0TAYZpTipBMNuJm
WA4iWKJPJ/2VY+SbYdwDCzlarCaZ6aPrp2UFkPVdef8NVN4cDeJWTPVdzPTgl8GT8rG5UCujQkYH
5gm5NMqYyeDGkC/F0jeoH4tHDaj5s65IoOQ3WBWVv7kfb6k7KnuUp1dGI0psuBZZySTMtzyop5ky
kwDPnXMkVNZADrO1X2D33kQ7yWEJNC0eUKa4rRxLPBPP0BjF26DDlnXcwyf6VtsmMC3yCSI0bl7d
9Mq3K6YgziBh+uZh48GBX5qEtN/EqR3RSQuuKVg81mmibRJBuSf56ux76wnJsq7afOxXeGamC1+S
99mYdOPcI6xfs9MsrmRLYv8cTzXDZm9nGfhM/NtMCzS5JXcf2AX0U24H3cvtqk3iSN4mYFrW66hf
SNeLUmvWOhSu4SQSog6lFwkWTkN3UUHUnSX/okJ+Kax2rUDCXDLYgthsPiFH7/+HOPRcA/dyRezw
DVyKe+d1Ag1KQ7iFLmpTAi4uUnZzM2DDANOa0lNVSuiqr+HJ1SlQYLGdcn9Ol1cEaoEDyg9FFp+r
xNhsPX4w7uw2G19IipH+5eHrrhmocoQO1gI7Ht5umYAt326qo3Ov89vZA0eEv+AxyprfErp80U6B
pNArhB025q7ExnO3qgNyLTjFoLoc/oCKVByHNnZTvbybDypTkxvCu8ga8kHmw8Ka2sUe86qZPmsv
pesPgtz8FDKdxt4e1pCYAmVP19xUCxvJaP089NJ25duK0oHouHd37dU3SxuCy+MZnaxqDtYDPkbc
mfRJdl5rteqRZkKL0TpS7jx6dUcB9QxAY4+0kq14eVsFy9Ni9pHdUUukyAoDdNE8TMGoXH9q3mn0
mqauNfnuBGzLXyg7pM7oiOYletwooDtgoxreeuaMru/b+pX943+up0PotFak9CC1//PR3xWQ03gx
j0LhfEMbYDs75j4FKL8bPcsYWvK/WQFIpI7P3hL0v5RK8aLdN4T3RFjFG5aQE6eWH/yk3pdIzb2r
aJWmx8s3jOdymE6Uo7wULeB58IPnyK28/2G8jm4sUyNAxXElsiW2HQvbUjdtpCde/tzbHwewRD/U
jUdKFGhl5TJp7wyYTKMFWUqeEqOpMg2zkjOIAupnt5EdOlQnJvMWe9BJShYtfmPheppWFvmqoSg6
8ghZcvlx8fB45dACw8zJpcNxRtbK9L9YbkcT7tuCVvfi4mc+KfA1YMYa2ne2hHQkakQfB1Dy0LaM
KHmdXX1NqNYbak9ZmccIvOr9ris4YSU316P9Me2NvGa8ikuJzXKF+CY7Twd8LA8MzP/MmFdUEwxm
GQrqFna1Va4LJbHFNLy3BoQZwGVVm/Wk4Z4kWVHwkyGBwk4SQBVpY68az7q4GkN1Zw1Px5ZDHQ4E
txE05BP1Afu2PL4xKqCQfsgXOlp4NIThGcQJ+LGHCVa7OivHvkA5F1oDzWKxPgukigHLANcQjNFY
45DYKTm8wBwxHvTrjKZzJ/mcN696xqiH8BLltbjPFoZ/fXMPnP3IiNr2lDsJWOa5M5IPS/smfLxB
kEM/DIAVA+bacY9TvcljZXR0WrZxd47NnxgEK42Ky1t6GBuhdHDC9CwrC+eqNEtZRlW41sXBLgXA
p+0iBl9cfA6xBaQL0s776vvUkS/mENraRwiVKxplrYbP7XPDUKbfZAhsdRMKq4J4EzUwzKVPPQDI
FoR8+WDzyyTY9M6Jiaypg+52zvllWKPljDKV48hKfZYTvaYHfMg7GAbFj6GrsnFKwnKnJBXNB74e
BWcWSwz86QACdWJo/f91pV3HzLt6Tt64Iw6kCNG2ggjmiIEImWFyahm2m6n/POuxiI6wwPiH/9pZ
3J+zt9pKu3B275kxFvbv8q5h0D9BnXMV6y7IGGrj+PwhNmlVod/+5p+cwgnZrhfmWwdOWaod0JU4
H1kdO6pKDYsG+TvQP7VMSoW0xDAP7xVirF/h1gQBEa0CwbVYNSszbgxqb2QcU7cPm/yFVXn0mT+m
TXNNr3IypnjPuIlSPhumHdpR0yog9yKqPkLIY4DISfwyOmqILfzTRdoOXGa4RvxgwflhDpLFOcXp
EdjYVxgAdho292X0uXe+C4rwjfvI5lx8+u81qBfE0zUK+WDklqVk3R+eXS3EUnvM0MFWUXScMuDT
kyKgnY5v9qd1vWC/QuUcp9YEoEXEkrTZCozBZ4vRU+B1ZrfyNeqFvPe0r8aawFt/rf21mzv1rTId
c8zb3w7Qbpk1J+ItG7kMs6/5u5M/YpnA3LUljspU1ujqP05lT2ilrigjcYSx1aoghw7+mxj+TPzX
5fbx4lcNy5sxgfayeINFdPm/lUN9W5gMEzKx8b1oEIBeEg3nEZoQYkvMu0R0xP7FyE5NFfsYM22l
Rs3+fwmTACtcfp49omxsqrzTNzNyiGFzysjdDnxEU1iBt8tX5JjCPVyPa+wwJi2WVqJsII4HWLXP
VMh+t6p1HiG1Cmm6u6nn/tIvvuvwVmmP94yYikbXah15m9ctQBC6eCBjoplU+nJTlbybuaZY4zaO
pNLx0+kyA1Wnci/ccRNN1dINB/bQNo9fa7PMoxTYKySds/xwnYviNAfPI5DDsLqSyePpYB4uxDOX
QwsDcH+YLkgz7Kca0cYWKNoeqgbr+bEFweERoR4w1bsd8gkmNVVv8i8g+/KqiqKDFnbhd/YNUvyJ
1fyLrP5dIUtwxzPKN+tkynhKXVTKcuhYSLnyZdjVO9SmdE609B22GJ22ol9tVARp4OYDEYok7p0Y
5BNhQ4sHoDsufNibGHy9WGjF1U8p9LnSNQOfNIARBgaj/RO5nzsiTHuUSPERR5QkUbBYUnDZaECR
Uq6ZqA3tpoCkbBh2z6XNg9WyDlXSB2I2OgNZHJ0VbuLHj0q4vhtpjbqLarVd1mrBDGF58HNZVaHt
zDPz1d/k1So/3+3ygNHY5rkTgV/P+yexdE5Rn+rr5IUrpwNAOurLGqbTdmyF0IEK2Vyemfa+TzvW
uash1qTEzj6LDsG/AwO9qPSmJxjTUO2Y8srGhRBOJctz7LOCGGcewcQkanlAeWYPUzcLDtzn3bjb
ddPnThWxhn3da3fgq00htTsI+vO5nOWpWVT2rMKg/FiIbt3hxTLDTRuBtXSMrtV80xlywIy2Bnh4
YcKHDoExgP9yCGG/aX0baqpFu31OAw0G53a50EFIEx9p2T6UXGhrnxukVuBxZQ9xyfqIqWZTBAU3
68IS4vC5dc2keHqFIiy3H02d4mXJGOqUcs5cAfWg5giSZSMQcBJBtAgT6GFEcKmKq3WINjnP6jhU
ZOi/9ikePOjHvIqYbXeArcX6rOct3fOvl8Bg2YXdADWO4uMbNDRoocWiF6jqoY3T4QHFYQWfxwAy
W57NGHp1bzapvhuzr74VkQD8hz/2N5mtCFkye3fvhTDuJ3J9jPjEt6YEuGr8BamiiJ0q78ej2vI3
V3A4SBRdsbbwJBXxZM5dLBbJpsoudC4prGioZtiB6Z+MHfWF+ieFjIdXqiA0A7dQ4KIKSGF1RffX
gulfIrq5O7z337l8IKnKtguBywPvbJaTVbm0BvHrJZ5pfLG5YuE4UkIYqdsz0mFwSNCZjmxR1wdp
WTbQriNP5+YarSpT9OCddIuL38SOUnBV3e6Rp7IbrK1KUUCiU5U6llSXm0b1OW5ZEBv9goV5InkD
P8DLL/dXjDgVWrBRNr2GdFLYiKBsOqGPOn+04HjauXL4y7Nxpr2pA8nOKCD5qSpHYD3EK1R5By5h
2ACERrjpJalyVUGF0dXCJslBu9Gozf2Milbji1Aq4GBRYcV9xDqhDE6cSeiwo+l7l53npbM6UdGo
ykBX3m5iCnyPVrQQRgljvjpBj65y9sPY8ZVLUUmUUXix04OmkLDsqcIYB3KFBehrc+ehT0+pIRSo
WVPpwIJgonvpRYznXQbdJrmcD2j+yQ1B/uO0xYyiVbxgOlNxjEOU8xD/SrYWEWQ3D1k/8diG9MBd
amVGo+kTdEzVkbMoaPbDpY2rgiCWiv5umFhB9V+f5pef/NjNKUWYMJnpUTFu8+3fhunyOvsPIm/w
34tTpNEDcwK0Uwb7KRj9cCFLoqG3CB8onhRElPaFoZuzWjN7pppgRY4pxbvkwYnIgPlQjWph2WmP
qlvg2xnrGBC66Vbndy/70IB3JaG7c9Zs/Pk3T5hDnhRkjpdg9eR5bVnevB1X954mIK7B7yoRYKz0
yxOluECcVJ387yIWdqOo2oecFfaPe11eej/vKnMIUhnZlksfFPQSB7GDOmJ6KXN54+oNxDJ7liS2
ttjYLWpoRRNGfIUv85VTkM/1UiqR38PSheHjtw5RYjINguBJhrZvbbPc4ooHgGAppTRImv9YXrj6
+/emBTtFU3buWmsSOIYae8YyO4UiIDtmZTGF2oJ2VIZCiBTpVqkq9GfPbiHINcsCcXWqd2pd/sjg
piETugCgpLwqertWKfH3R1yx2h6hsoUZl9pD39Vh/V7Xp9pci0v/2FuViSumwAmsFk/6j1nJMcEz
VMkNV8zM6OXETOYyxb9FtbcK/nbAU1GoMJhGxL1Q9TYSbwlFvc1jrbuYRzQ3l+D1Rn1fysDrdiiT
gAnZTiZ4SV/WORxIN0MhoAM2imlGQ3fHzHS8Cqq+//J5vA6IPMccUviHt3lymhz+Zt+b/0ru2eHL
addmfPqNLITfphg0tlRfm+dOYs/oEUSEvc3yYhKr/GTP40AVICchbQnj545e6H0ECRq5gXWrWZyt
H5eO1ka7wz01uOZMm+XFIID9LzwB/rj8mMWBAzCdSTrmS41pXq4sgz6FmCHNQodS5LpK/iiaXCdy
0cg+0jhPhjYj66vLTxm1WV66DTlZl7eqrcUR5Y5GJwfcNzu3rbZGgM/G2t45nlk2T8aivuHXoZqb
stdk0szxv5Gv8iminl+RnZycmijllLXBGSW5hSB34nymnyljyYgwh5eky/SVa9X11TPWgWUkdh+2
ZlSdGgNMu0OVuiqEWn9PpgOKLhbIo1+S8Dsp5EUCSx8b3CGbBrM3YcpcyxgReubEKjWkL5BUxqho
mPbZvWiCoR5Jo4m65KbbVaN5u/pW7BMyBLsDrt3p2boyWZkniYYYY6ySAvSDiSq1wbtsOB0ariM4
rn9FF1rtUUu7Qnyp/WCUvSMItQLpdecw5FySFD6kdWjyA8vfAysD1lCI67Namco8v0/fMdHfbVt+
3CiRb7TvnMmHmFRU/qB2s6zY06FBhfRrXja3pi0seXbjOQfrPLwSvyghX3m9z1z1S9cmeD+UWgzF
9xEvbesxD/NJnZHuJzN9utph1kfQwTstECJ++B5WOe5615qF5LuIw0iFGN6ag4u2YQXW+LjMYtsj
pnREk2p9UVJ6T7FhlItB7l7BVFwUwRHkjXCqoUcl0liY91QkrLFLMjsaX+i5HvkBRmRUcWwiYx8I
tRM1COZtafYPkjiNDxdUeLbH4aJdKjDdVvHbgeRtqLhO6z2tD7/hX8SwBEXA7ayNYc2ebc6xGQ4s
IFzLDOFkyLtcmNK5H0qUXaLpWEza8CH0+egvAd7a5yugHX6p8fL2OOQXT0wc1lW0USUlA4Z8Hulu
Z3n+igobc82iGBhkigy+UkM63p9i3wbRrv2WhNtKmlXmHeo9KSkV/xQbWQY1rFWA0UZwf/MIhit+
tD/6/H0wD466P9nEn/u9WJg7nDVOWGD3/cMnYxjfSpumY1zGXDC4b3xQLUjBL33fGRQ9U1tUBi8q
RVey8XW5CraVxnOLwltDNEIw0QRAlmbkDddW8s+xQqDOyzUpgIOkDQfWi38AKzPw6y7UXO5va62b
rvZwcL0lDuwtPpgfAW9iSlD7U5PpqEu0pV0jPDNNVZfwn4Mimcq9XI7N/sUrJFTA1V6PbpRVr//X
/w3K35HS6NrTZq0R660NiS3HnkeaLupKapEmgUru+qeXvTJM13U9wfi7DenAhleDAUSbdcyI/sCr
xcoNZ+e/GOO+MChfoDdQg5W3wrQX4rIhpKOOhwsWXfynTSFL0ULkirNhjXkah84C9CxEbrg/lAhT
lvDccrfGkWwOszXCRrREA3fWzR2eS4wrtznUW/a9XS0eGzS4RntavI2PCQtB3iFCAzzfJdWLvaIU
EXhM9J8DyHi+fVBLcSxb9NHdHf5FD1bKKsM1BmPhi927ij2LxXkrReMq6IROThoEp/BKgPBGlRUr
qV2ZkgtEWwT0Eb/yMtSvnHLIiypr3f2yqvOU8rnV5G7Yb+ByIG92YdOnk5dIzj9Ck2uy1/IOtXZG
twWq3XDXcN7pL6meQMgXwyPo+qURawtcXODldtjUgVyxWQFi4IUkRdGgwmduRBU3WB5qynYXlu9z
duvFxd24u1xWlmyYopvaxeq/HxhZSkkzgVAjFO7Q7eUtV1JZu9ircEFoRRNKgNeIz2VDDGNgAud5
WX24ZGK5qMSw3iadlhjJAc+i43O1tVpcyKkp71vebM/OQ01/i8tSKJHiurv2fKPkoM3f7S5G2inx
3lNMABNk2cssw82rKqmdqJio94FCBMdzFHh/9ZszdX65b5VfhzmjsYbtrQ0LsoqiEQRhRrH67v8c
envBlHKefBQKogZPmvMn0lLLuJyki9PhQkGLR460/8l8gF4EpZJjpHK/fJ7CKwDvofcDJLJ93PQt
eHdWuB5uD/Zn3v2w9DsWIOdLfowHk6feELnJGl7+OaDektwYdtzk+41eRTbRqdKHrtz3BGiDl7+I
/ZTayjoWDj1AxEaWnLGK2UWamKoHE1yWm4z4TpQPUT5iYjyVU//GV7GeujkYlfXI5xt3SKOw/nSl
ctPVm/BzXiTbgS83Nn1bf/GT8ZVcdCSzSksJcylQ1VbuPX9fPf0E8w9W6kcNGrNDjyY591dEpcU9
WZ8d+1Zs3HGh+4ej7n4bDOh/CUWrVMSOj5oGSL5rh5APsY618B5EdclEHdsXGj9CGZnujIcZn86b
j3Hg+5eU+dI3bf7NeBu5KhiiJ0XSqAdiLpVJh7RFI+2J3yZLyvKSh03iiMubjcdAzdylk0sJMud1
Eyk1d/ScK4Wal7bazxwVBv5ttWA2JvJLjQTqkvPqXmlWilkt21/LNXJSpI1g1WcP4lqSl72asW1V
Ja49FzKURKls46N9FXvpZazkunK1xyxqn2hr3WGuvI7gWQ72R6QCcg6LrNQwPT1BTrko5/2cqQfk
yf3X7jJaYirtd9umPGfKGx06rSF5YlrJJMC9Gg7j/qdItXnFLf9C0eCjEeDP6J09zR8pz7cYEssy
0f4tRICAPt28CASfEH5RpXSBqJg0RKifPK41b72NHw2Wxv56Zl4XIFo5ee6TdmHeXpqoxq3ALhkj
4kvq5tHWSrlqYxkaW6xZz7+eNClrWVyNpMSImtwl5hrz1UfWyF8QB8RCLzY3ZBt9DehVZLd0nqpT
4RkOeLN744or7Lu4xUhYNvE6kUJVFqZxPh3tzIISk1X8rEd5fh4Fkk/F09rUT3iIt/Mu1XmI8O8s
qsjzOFwzhnywnILl5YMXqvyxUEYKC1LYJKsAzBdIGBRH5rd+P1YQ2vK9SrvLUGDUFTs1pHj/iVGk
uI8yw34CtUiX9vR34xj/2OcjE5rJdyFh4hUxAUdRp5lqi3+aU1jRNRNLwkNH/UdTDii5arEIGRs8
EmVNo+xNSfah/s1+WIC0ha4hW19c8NHTHnUDyXIgcjOSdiSAlAgGbvZcTpP65whVsmgYCkaVWNQ+
VMm0vYWuJt3PL7L6BgMwPgXJwGai9RXihBYZ2C9ZU0VSynVnjE+xLFC7nmcxrL2PdYg985qbPxjn
GccPjy48C3mh9EtBaFjcTAypjQuYgF0Oun//jR+RymNuxtSnguhOSUykhlK9pSjPeKGD0yi6+Pu1
L4tD9zcFNdlPI/il9JmjWCnSCW56ZN+VbmYX6nsCkXJwZkHwnRTZDRaWhAbII2GvuFcJVSRBaFmU
B/x/r9ncu1qKddQo0QWwXPHDMtgPsB/ejXEr3TBgmYs8HzjwX07YLEi2B6BFWJNhHF9vBBOry5IN
BA5SIHuuO3LIrFbmPdxTBezfrQIgXvOM+jGPumhtUdyUsJtvBvclodOmSr9S0GnEZqpPylUaXJOp
GLASPOQXNt7KBqf98qnNF40pCoonwqzDCJOte+wiAcnM46/qxQLgUoSyIEHcv/4O1gzhnxWlFssS
4orpN44JyibTuDpiCdzR7ardI+fXr2fQXfMytyNEHfCA7XakHtcEAL8+kP/yU1HIyPr9V2R42n27
XG+j6OcSaeWnz2G+cEWd3+bdy34U8pkil0KAst11vWfAchN6Q+IYgFbAvaPhuZChtsLuNp+eApRe
RmRg+m+k0SHFSYyoV7TDQTIbfAh3w0gzDOPWkdd+NOFbPe8w+ULSKlh3rx8JMSf4fl0a72dz/Cut
8gFGDIVGjC3KL4zPtQBj3hupsw4LByDSPiGmGVXOU7ugMPENC1NxHDYkKqODgXAr35e3YazR3/N5
Q/PmiUxNIiUPAxe7OKytJYrTvjQQcTAZ4ljZBBQJPcjW/TGp4A7SMcSlHue1igmNzdpTX0epCcH+
w/RKfeGKMalt5xk+zmkbGu6euUc6bQe7hnjDWrocjwansuZ/colYvnRbJomaASMCgy5lUdkpap3r
Dinfv/TQR4cpedPssFjAINetSq9O0yerM2GeFTvY3v7NbhZ7AvoN2BOgdHMTxUToRy1H9xED7I0c
y5a0dApfuw5GnbCJLHR4oxeEsTSLKiRZq/+Mt4UoOVRlacGf+STBQDk6oHRCCcpaf8qLCX8yn84z
XewHOaiVZdm6HocFLYNrQlhxAHAJisDG0cajxJT+pl4OlyojGQuKdAiFVxAXmCrSgdj9jjLo8aki
3JrNa8LHOHzkk95bbKcayQpZI7NY1dyLaW1CCsjZ00wRr2T58SZ/2P4uV0SWh9Mvx59ydJQkVnb9
/d7s1CjTXyV97celY4hEmBB1ugJFs4j1zSa0R9jup4/7kvGhvGd9+mAyHAN9v4bKr3046OcBfrmd
GMdkw3dTB2S4YKsA4hOh0DJ1dk70TwN0psBH554KfisaKFey921kfa0lpPRosCVqib+viPXEjofv
7F1p1ma8HHfQ7XZ6L/Tzv0DDMbLAC74+I7IhZqKGTgaybOZnQe9AhmoUfepgAZfet5DGUfaGZCKg
wZJz4N6b17x0hOOAxJU2eOrAiamyjBa0Z8V53LeibjPmEwDqalRdsqHsHbkWg5a7O7nf5o02XCnQ
ZRvuItPs/GoK4raOJGT9dq0HHZDRctUk07kGb5hww0PwkGM6CNrzujuD/csu3v9J9Gl4YV2SnM1D
lf32N0HU82Ii/uLfuBj4jBLOThUHSl2ML2LmOjKlwu9w6vJ9jSvID6r0I7RmWIFGDIeT6jqWg7bS
OpsA9HW5N+fkFZG/PchbMmAqspq8VM8bbhyoyqMSl7vdnPvBbioOveTjHWDifQg8WwS4H8rL3EpY
sQAEnLNf2rciUcPxOf2z8G8zaaaKnsK6OJq8UcLqPfn/ueVqLr2WjJhljcj0jfKspnFexiCNROuZ
z6DtbOWfhPYgfjt1qIwifAlRfUCfQOrfGQy2jHnEzcCqF+APss6AaAiEPsbcNVT7zWR22qYWeWZx
Uwvm7DqOwMwL2FhUmu25ZrXf1Dozah2F6WZOhVzFzUXHoljd1VF9SWdzgCUjJhqieYian7u24zUm
cTsiVCeLH5B232P1b0dznM4Jvjc1KkRNznnAdvHwcu0bZWGQeVSzEkoSzTs7/p5zQqwpUD0NuFsu
VSzMq43lLuOdSQ5zKOEgeVkAeEKLZL7qmLLVYqWF1QjmcU5p0jKhqLovZtwf552sObvDXh2U3D1l
lWEwuT3PuIdPtucmAOT/O4AOqJzUyI942wg/s8/vu1Tdvo8cse1scXlBTLfLbi/COnAqgpEr8kYc
22fdg7IKCf/MGn/MLsQ0ejy2V0aAXFwuMzxlov7V9x3KHqebM8d2S4PiNFE8J/qwlbs8et7f3HZ+
TZuUIyaRMFr8fXddZSQGJKrN6SkAdXc6GX/owv04oOQ/Se2KP30Xm4J2K71MReZOmUAT3fwAlpYe
zE4n5o/1B1BBpyXWaB+nbW1kVasdSxRqam3gyxWWLQYZNnr6qpNODmZjpLyeRmkBU3k/URDwK9b/
r1tYpbLdiVra+WnQ3V5It1cd4lVvC3TlCMLgHumT0fYxqq7e3LKCrGlTL7qmn0VqkaNPUE/ZK4+b
k6/JhY18ZM+95Bb7TsQi/qWLsKJ/WQBtpK5Pt3qvmwUNQEnT4OduRlEYP62FHATY2s2S/D6LV+0a
ReG5U0mWbtCwoU4kc9FTD++jYFSm9cRbvw3K+t8Dh2pk0iinJZP2JOje7YEPDcwJ3RkeVLG0LUeW
M6jCNU+enI29Yh4Yv+SpemuUCw8Mb/m//HW4xLpja5gBVeWP8D9noVYFmoQ57zfvChEbuOyPr5nm
1Q9gnDcWUH8coaDJWNl969hXBjjwA7oDSaz87wL0g3xUnvg6EDRl+oJIvZ07thn7EdtpKPMJNK8f
XkbrSgNVPvjY1ueJmDvciV8s4o4PATZn6CHkdVuknzPYH/OhFrpvAYS8mSYkP5NWEC+UZwGsGFK3
opah6wojDFfeNwFXkiSOfmHWpgaDxuB0WETBAwfSt086RpgLWbAj7qxScqMGiIgVrB5h5zaROGqx
tQ43XStLOQ5YgmTEkHplb+flAqnbkvb/8z5I7NjdeTny/CX+ILGJVHSfDFjk/jqDYE8+/uj5U64k
wDWAKWfALpNgXmhxuHmz0GUzsy7hXH398QNTu60uNRoN6+7V+4iidjC0Qvtm3FhtdkANd1+GbVO4
Ome6Y9efsE5hPknEzWutPtoYwk8FGOtBQlCoGWPqIanQU1Hs2A+YKcAjRhissJsQvZqocgnPxvAT
zYIkn/sc/iA+XCFrX9swhxWBDAVhixW2813RNTWlwyI2drzVHoWOjtB2VCKgYY6soAK4Aqs3Xza7
zLgXvu6goQxksb0/PWkilNhJqTw3yd8nIMZSVmQsHRmCW6gQCTf09OsvEOlCtq49MqiwXkPoZ2oL
HC0DvHC3+gDPVPi9xOGd4rpCa/CCYdghg6MAunfMhQyeeRqL1j36LAobZP/MKgU48cNmCAff1/4n
7jX3XlRBARMcuM/OLQ/z/Irv+PHNMFiph4t66OyelgCspdk3FhYBzQfQPlFuOjJ1/ln6mU2B3gv5
Ze2RatanQ4VhL2KHCk9B+B62UHnrk32Y5lNn8GCZwkEjcDXtcR6pmZGIlBzOSFiXLVYOG4cRUw3S
OAON5JhKZcW7UDx0KkwT7DayZ3Fl8+zr4RPEDIeSPe0eF1JgtgzoQPHtJGq5fmM/H8h/fK3hg5H0
Akouts1PgzJ7sfms8+ELkHeXFqCeZmBjN1U7ujqrYL6/RLGdKOIjFA1k80ehlq9z4gzJYmgw5she
m9QbFcO4/6RZbNaWo8Ug5O7hMMgFxELsghDEPTHgQywSFI/dUkn5rE/+b8KYO0KrYTuufUGn/jW0
WlhAKP0uwpWygBlVZK+7Ygjfe+uIsZUFINrxodWU0vyP6yDejGjGJ+GpCQ9aqKPjfsBQoHtwh5pl
FMoPn2RDfYyIFyayT3rdNRlCS4i4Fa/NdnfVAWpVGzZnVNa3l6UsF3UeFAmj6hOlleS+wKqiWe05
krlDC3b5igtxAp9/aidBYktu5agriea5U2fZXGAQgyJfZ00Lmy1tB9KYKiDt550nkRj9L4zu7dfZ
tMzM+qZCzENsJMP2Qn2zAdaM4oS7eULBAxUcgAoaej3k4WPioktmqm9LfGg8uzjGNompm6dyyPfU
sPdabDYl9jAo2MN69Ly3Md8OtEZfI2uwgIbs4jU2APB4o3SxoU3fx2L3tOBKPArVJMICXN06gy23
d9l7+PVuCtyX2ncU+0zdu7MQrEmM7aJjENL+Jg+ZyDh+2p5EVWogk9L0ZG84y4HqaqLDeOVqHI3/
+7QrVvGe7EaDRgaXuWoX/If2Qqr9ukQ9u/Mw5gx5KMorsQIXf+1iamA8WXpiqgCdxnOtVoqf4j6v
BXCCQSGDSXZfizTroS0xUsoQFkOqz8fEFDu2uG1iWi2x/trHhcrDTGaHPAwyIDNjQCcekEwSrSxD
y4iVUVGowLZBrA4PRGqlscJ08svtZecZSK5tPvnNZid3OBpNm3+8C3s/5cbdlukexSwoIAgrZbLT
IkKR38ZrQPaFVFNSXISAsElrhhDPDU9Ekl5tNJqwkT5ErR3fw0EZ2J073k3jdXiUwLdECfhnlrbu
xF2ll30SP3O9sMHITrV29Pcu4stMnQFGo7dwgx6Lo3lBbcCE9/1uJ90Zj6ehm8lyj4mefxIREu+e
VY1tjEctrhDwDbuiIAnro5pN9ZVCNQ8C0JvFdPX2T1LIxphhDtyfNMEASYnaq07sn6/nwrrLehId
kFuHXZEGZp2bswQfkDh61MXV+WRGHbveQn44Se1YKdLd92CzwgjqowancYdAVcePvpS4l4p+VQ+W
IaAhIA0sokJYKBGx2U6AdI8RFG8wNpPPDOpVlC1G527VEKQzcoveRBOUuL4bZCOkaQILQVgCXklS
4UqQTvT6xtlvVH54e/d0mRo1knNGl+B2RgFZiXISyqOqCGGQft6tO1OMFBSCp0tCYEtGZdYy3IH6
54WK9bY1ySTOY3/8zV3tcgwE1MLM+9ZXX3Q6xN9BZwdLoA0Vun0GwgnquLmqdjR3z0R2KWvpNrJQ
4zd3asD4C3s1+ZbMzpo2ENobsZN//RSNHCdZ96F2skQdJeXkat5n0aal1FoYgCCiWSppoO4fo/Lp
Re/lpOly5OdycrXp80ti4GOkvDU0dkYKu+EO+/TKvDJ5EiQLo90G5bGpqaOEXVJ4L97YZrJHqzIu
jj4/erAdhVs8zZRu31YXEUq7HOaJBcscZh5rnZILD9fCeijW11eM1/tbFoUYkwGaodG+5uFHRNcN
WqeVjQW0zw8yUKL4dATglaurE8KO3KNFnCjV4vIWAz4Sas0d8h5rwujrF4k5xxwpubME098wm77v
it+cAn5oWfNac0hMw6fqIMRWvEJoFv8Em9dIZ6g3pgO62UkB8eNzCO8w7DdlJ8r3e+ugsIEEPRoi
bEcaLr4ap1kwicl14a6r/cRQM5M4OLmrm9NLYF+g7OggGnGHdC/uxPLlJuvhUWnNbH5DjaDppiJw
2hjCe+nnVB5kUExq5IdiZCexMMDp24soA7vRXuRtdOg2nhID1vHZLBLW3A2LvTkHG8XZ+cDDTUjp
kxCC5W/+Xlk5jV+OGtDK4XjilXhJZcZzhSs3vX61G4hJpDaBn/wIgjgNE6x1QbDhNkgno64v1qyp
aLZVOm6SJimj6zWQpAsSk+cV+TfHjVG3fawmI+bfc5HWM1jvIAJ4zsWwZUPX4Uaj4r5jemEKFaG0
oFpJAL1KYoaANxMXVQTWSKEkt6rlg45NaV8znUoUZToodIDOcBl1v4zaH2MxJ43ue3PycecpyloZ
Kmd7v0W7mkZAWkpfURnuniUc+RrPmwNYFpMFltQrKeFDHoe96KvGfipP/eqHf/wu63TcvDqyNLJ9
8qihq7u4zb0fl9nECJxbyn8dspEbW8g2vSzlORXq71MTiR1JMPD27x44li3Z8AcSW2XXmBTpPK69
mB7dmqiVds3Xgaqdisz483nCSaAsjrUFoSqvIAr8RveBVnlblMEy+tt+IeUYD1Xut4K16IhO0ed6
4KHSHNUgjrLXbxAC9dKxCbTKBCRCjYu0/u8bSJTSKk1VX5wH4aleZnZVqQvuHiniY3Djxxk/e9FQ
k1ifvgUo2K6mnSlyl3Zb+33Kvl+X3RavVOIrpqRqMOzYBu+9684/YRaRUtdFOmJxguB2wI3S1vkA
+pJnXTDRaOjnw7UQ7pE9xmHgg8JEstGnEtcHDZg1S5RkGTVOxLDExhE1MZG0HdcGW2v7aCkTK4Tm
LyeDcQ2r8EPC4mDGRLrQFQc2qXba95GcJUHdg0pJ9dEyBgKMQirQV7RNUrUUslSTHEz9u31+qsqM
ijA713IccV+t2L5qspKylAPjQwf2d15bccHTk8j8Pgm9b5hb6g60+Ovuklm4/fIx5KDtc5E50Hdh
0Qh9n7WAVjc8UHbCn7pakOwDevPy/tR6qg29wVm5oemugJeTsHjmNdJTg3NwsWA8sdYP0OcTlLQY
98V//NDL/6NWSl6Sv3d+xKQS0rgkq2x3F0L81QFdnbwE1xUKuKp1X0NEc3nZkXK814nAsZE0khsh
N5XgJibkCIJqtkD0OnA/VVOGS6qg3AmzeGdq4MzVwrzk2PhEC7V8oahuqnCk5oWE1+muzdvSB/iM
58EcURufBF/7TVcRx/Neg5OpJ4g6/xqUUaZlshk+pvYgfsjL2iWNFhFDP4YfZXQeA+zsPrKG/NAs
0k0BDB+gd/vin/ipm96s0+c+EyKFIwZ+CsHUHhBm7ABDxNgVrAlTtB2nygbQsVFMqS6l6qHiPBYN
seCOZoxn8QxpdtxT2PcyYpZHkclQ6zUX7yl/TchHrst7Jtz8XJS9f8Gp+tyNJc3txji1P1Xwc7Wq
/2imkmQHNzokjLwajYcuAfvrGdhsQWyRTsAJwBc9N5IlIfnchftIq+ZM37g71RKTLumMLPX/WOYG
CRpZ0K1Wze3AstShrGQC7jJO5AOWskKXHKn0LboqsmvOleMxu7iytUkkuQTN0c+R8kYvJGwYF0xN
puySz6ySDCLhLjQPYGHVnG4szmRzEl4GlAxGm4RL1g5jiMw8JySi+IC3MRAqk9W4yFu4jD5gzU0p
pKfctgg0KZlq/UqmhbtHvaTY3ak87fAxAo1oEZT1RRFh35u+lg7mC3eCUXoHWeR3zRa+qk/pcYvW
CdCelB7fICvc3tzeGymv9XcgU4Tb+/GC5smKFLTUybmstvAXk6LFtJWpoSEUz5pfdLlXgjCaqMY5
9k3+z6dUdmxECyKgMJQ242SUJGeo7gpUf5TRsaIslMSvV91fracZvidjKVsDAKWA6JTmHh1lguet
othOfOf8JFgHwbn+vFeCn26brjtB5lt4e5jvI8C/A+66Oq15jfX0ekWuzvuhB/i4199npPABIz76
SAI+UsJfcbSG+fjT8P9Rt47K++p4Qfa8ffmiXk6IsTmNc2MDFk9pXFUUcP61mj+3E5bR3BKfDI3k
I4hczbNsWUsqcR4u7nK4TExS3ULytNEqHftl7erQDNQx9jd+/e9OZXNfzMrqzkLJjDcmMvP69vKR
MfRJP243MgzCj3t/1dFl9TqJjide9gBkBjjYFJUhgh/ASnNkQiUT8muPB5trpz5ELU8bPHLJZeUd
NL7R0ZGL/6WIsBH+Lh9Wppq5V/+Xnh83HvUZuEvqloXD3EtEwu6KyAn4UPRU/dkSrcDoHTf2kfNj
KKkB/0mhWfCNm6VXTAy6nSxBrL184UEnJifHRUPwdpKoe7oEgdmC3jWGB2bmS2GRqLaiPKLhm11p
ptzjRmhYuRj5PIIucNxsyLCYFlwsNWXjJ2fVxM9j85viP5wqlVkhh5AJ0DYSPGKnp23yM8yvO8C/
aUW4oDrXIeQTL2EA1ypQzZHpY67Mb2mnM4m69j/KOkbIa97gprspW4CjiPo/as9Px5vcJb6Run/m
TpDa9kmqWa1/MyDBkqV14Yl9xMTbjJ+vYOvlKuHolI3jRr6brKA730xaJjJuBwdv865+5z3/6nSC
NsHGdfyTH1cYMfU/2dU60oV6QQxu6ro+YKP3SSsELRt88bEiG6QU9PU157KmA1bMMBmoPO886nxa
JUB5io7vl6xWic2Ggo3DIzNw43ylV0y7PsNUFTfalt/W12QAtz3WchWX6IvelbsKuRrlGYnwQ9tp
BA4RlDNFz2jOn9Ju3nMXfAeSPnw7E23SGOFyAA3mpZkguJ4jYaAIR7M1vaR2hKP6l8JbpjxCRErJ
dY7VKSJEle6ktE/zyvGYA63BjjMn6b5mYS3SJL0D8az7UimRr3QRF5lZVL0lgu8xOFgqRQnhZ4rs
C8f6MEynETt0DbvNOOquF7/rwhb6Hm0Irg2T17trmAfkojPnATjs0V8KhIo/klFRQXr/t54Plhlg
gQL9ASeOCuNwC2PkCxMDEwW/mrbrXQqS8XFIVQG5jTgAmVR6W/K1UrVHQDfnnIzMayhLX9oBWQkL
REIZbYgWV+UglpOm6kbYnWtmRmvdk8ZyfYPtpoFrjaevQjrfn6h6/vOE72zgKvkEolY1xhy1yblq
EhJ66vBvKdlZuUXRTqi9vI4YhCeuYR6paspu79/1XgU07qhpZfDR9FCIM+0ts56xPs8kovZhGtkz
c4YtCIhisCvyuPMERfm+wUhdhkae5UbH8RZEggj4fKZJW/MdGIlZFrv+CIFRwavDpODNKiCOABjn
LmUDJd5gY21SQhVTDjbF6+Gq1v0DsRoZkeWuyg6TlnowMTtzaKHnJRTILQnlNEIsDMlE2vUkRh2H
ZMPefGwhkYeuoCiMF5vvdDtoHhKbG9ih+NhzT7ZKNqR4bECKagxOj3s9i+QKfth6pK3OQ2L+12sg
RGSwaIQeI9CAyHNrrJA6FjTch7IVG+kOAYHa3ehOr7g5tQiTuToYqujDE95tR/G/Nzds+TLoHZQ+
Kbj/ByQY631bgMGfcXJAfvmRkNn8cQ4iOvdpPRCPpLjEn+hcecckuerLRKUr8T5e6kPLB8GVmnAj
jNVJxP7X5Z2xFJKvZq0at/6sSeDTvB6Z+0PwArq/AtZSZnH6rwjXahjdXK7/+bwP/SvR9bqw4o43
UOZsd43KSaFYuw07Jlva9Zn4cLf3eLV72iCRkcxM9JDz9ocx+6OnRUQXVOlHCBZH5PET1slAjjdm
oeAYcct4gWOFDAdXeysPcj6XhkYm+G0W3/76j2LeT03Z1ohoPr/4koqbeG2LQqWWN0DBh8eDfsg2
uRhgWbN0icdPPM6vdSt74JtduXC9Zz5rEjF/24NSYJ9c/9oUozKKKgjjLlUdvjgw+SBgsYIuthCq
QQijrxxd4Q7kSoiOcj2rBRiMsqS85t0tAjuR5OaIJsio8gQFTLOuMzhALOUyVs91EmSxcxHlyyHY
Ljukb89JarSrmqv7pBh0jgA/P0JEmO3IvP+J23pgt/YNPFvC3pvetN7ORz3cMwk5xrclJSPkzjNv
qhFgA0XhyrETwLXdwDcgrYwa/iWjKco1lL6Srgxiydn+SssC9WGCnTAi0tqnV1tn/n/qA456HwnM
4690VZTPEVTz/eVdb6qs42159XypIAru3pO9dcVPq8Jdbp4AVu8jnzpO3JuO1RuyyzQ5vLnLHP+H
VHZwdAMdWyr/geM2nMX7UytrCTcn5JSQ4gUNFMrSZ+IWPZlA/sdRh0Zk8CoGekXkTFc+sFMOxZzT
p/PGy5ka+AnOPeTK59CO376FfDjF7Sfgwt1kFHXnBUGdpvLCHkirPhc77sDvn+d9gFeN0+919R+7
Sk3i51kax9Jl6YP3nABGAEbK9yB8fD4eW5Ud4TkmyT7Zl2QNXQf5bn5KNE387guJZrHmCcTlwfk0
dPIpos008fVFrRENFH47Hgws7O++gYAb1PmjfOWIWEpwt7Krh432FNUlFThwgjh6zG7GekNk1gOR
q6TnL2OEn5nXnRHr4uWVSGM5aTu5yS3eOPccS5FkFKrpIHfSLIQDhu1UaglOsE0CYqsEbY3yobf3
9jmMXxZeTk8AayVafp6/4x+t4Z0uWXBlYyXTfa4yQguS24GSrL+G/2kZ95BKdq/gn3J5I5ybDlxZ
DBEvWqjP3udQCOTn/p3OMoZnx1HVnLCQNZaDgSn4Ttjc18HmntVzKDY5CnCBHCNbbe0hQw7JqHno
8c0CuUSiayksTonx6fUdKrFDVfR03cRxobcA6K71VDxNVyuyO6yKJhWcCwiAfziUr4LSOeUXg0As
UmGY50xsFTYReP7/upnbrJ0CWVOs52BzJ6TRlGNVcM7a5SJQEtS3ho8LDPCQ6A9PWWz0WMy3paJy
s2ALO/EXhNdeXDHahxuRQd+WlfB0NVLbYh+tIPpApB1vTVDytouGZqM7alVOss4rs4TkTwx8Oqz5
l9CEbc0XcSpx75ZvSlWRST4Q72ZFBG/DxXHx5u5XXj8TML5Ovphjy2Pymc9Rh1dRt6kcwZBklCAQ
pfiJ190WhHnPtcHUBtOhbBnScZrtsTl4L8rr3Uxz2dCLrHfNVQOSE5PhtGXUz8R1Fsv1cIv7xrpr
MlSzv971uLwjjCCR/BDRybrxUCZmnOhxFR+5vrNvDrnw88Vsm3F4BFp+B2A9Eo+y4KdG/+NqjQc4
i0pDJ6WU/v4Z1qqRV1FUA9yKVzbLcuW8dUwTP5nb5FlhfLDIqj1f3+QBSwElkJwR4C4oomxOFt9K
bcTUcn9xRvPlpQKRB+NOXM1h/09aRNO+pLJ2j3HiqjMQC20dTkshV52MmFlwsQd9c4kpRZT5a/CR
TDTFFOdjBRTQ3DmJxtlFMj8xUDWs0rRS+DoIB1JON7YEtqWjiUnDOoa5S1HxGyQUVrNTgttl+v+f
VPkVJzDf7r26jD7aawIalH2PJHnE7uzx8ZHUuyesO/KGUDpm9BvN3NtxAkkEqqGTKvEaxSZrynno
gJNEz2WJpYxX1C7hGyvDA9P2Ow2+c/dNa4p44Fo1PDosUT7vrlCVRR7g97bW8M5EZqIiPpGP5kZL
TcmzVtZGYw3jsipmo4vmIYmKWdUpN/vZnR4vdTvqtZxnxaw6MIcI4j/j1gatbvSr1N92bFxmNspG
b3HUYWiB6XrHZY0rnt9J6tEcd8kXyhIxYiSIe9r+R7DDTHzSuujQXy7rKwaHddPvNXYiANzhDcZ3
6BYdiaC1E2qkA73a9b+EJ3skjeKVga2r2vn6fUnQueYLie1kZxJkEly63vQ5f8gc7NtoxcV2qKLl
EDnFEce3ozkg5Bb65tb5tS9/tFvV50JO3G+rU60HcXmlfXPLgYLL32Eb/+WCwKulUEu2kln7GxEK
DRAIs5oACx+Kkq6suGC41rih69sd/UAsiOcqZIb5r+jzlVUL6sQGz33HCBMjfAj35c+kCyIJ4ZCX
RL8GYrv+JA01xWTeT1iMcZPrVsByYyTLTd/hgHVDiyV/AgE05PAR4BzBeL004ZgoDivayfuToGiF
SCucvA1n+W+F7qBJlD3vFoM+nfaeGHtrsCpCRCsXmvpmTX7sL/NdEuf9ZMI2jNReRXpYncxonicz
Gr34yHg8gZGIgvZKcYuzFjKmWNtR+hZI4WgZRDIzg2QPGb2k4hfwkQQwcI0/T/CM67uKLiKYddTS
Njlvci3Qa72TOtT3fDsgKIuQCqg1xYSxF+lrI92oAb8u40B4f0ALai4ig815PGMns2ZATtJ+L9vy
3jl4fNdMI2qaS35tldEtKYCRXL1F0dgDD+PnpyGSZ6zYeTDcADnHe3xcqwYdMC/b8b85VCTX22Hn
bAhyzZRe6rz+wgs4MAZmTpU+gVf5gwlBR1dO02yBXqCgW14IriX+YQKNOa8DXB3Kralsqm2RZPs/
0cuABgEcyMda14bcPUmbZMMqBuCG6a+2KWIPYXsoHu7qLIBOwiCG4We0gZftF+JzWKKEMklfeJNh
wrsOL1jPAR6yqiJdyAwRpIB+Lk5ijWAOkWExIKEfalQuzzho34aLIyJlYPqvmT0Pbbr46hNMUBhD
2gMIPSMX+Zq4p3pNiBBTVql9R8ZjtfXm/3Vh/BAT/TOt1Z4q+I0dfImVXf7siGAj8J3/jICck+zj
x0Y2zz6WFkDmZ8lNij6xFj3MRtlZuXFiEUBFf2ACn+1vBm7a5aBQCo5pfIFK+/ksxP0rqgL2AkJj
/KFdpxKxtvAPUCeeQ6NtnIaVVRpsdK9UFhKJEUV8Y+LrzblW5C6yhjqvpgstzrg9E4SmBKFeHWr+
cBhn9m6IHxkVo+qKuk5XFIOFiksP95KwsFT2/y5Ew6nYUt8YjVZFz/q+2zZZmVYWVj5HKpH74pvn
d3rcFYiXq3T+gnU8pE5A5wWgUxw5NcfhbnMBl3bw2tXKoVfZnWyp2zWwz9UwsjSNleE96ua7lGWe
XTfXGnNoUvlW+ncBfqZvAC0L7WXGMO4eGSO4N4M3GCBInpgQn3RVkyCRDHVWY4jiRmcjN5P+/cTb
5jNvxfECU6YVJaczHTA6BqfMvq2wuSGw2CFJ48fTJ49OjQhRBXHERL1tcQJJTA5f6BIJCodUcU7R
jNhZPRAUAccaonvbBpL4+llIJv9khConvGsYcf3emAKwibESQWUczqEWvP8tEJvdXwDUJQqC1Slm
oQoEPTK8xGcanEaioRjZIdAraQk9V8dveT9ctEEx9Y4P0W2c2x4Pj2pL0bfA1n4LPLYMPggjv8R7
jfQUMj87cMmszi2c0bmtriy67QwE1uD0PQ9UqOoYzs8U/d8SOlBHg2cXV1vRXjDPCmTE0why4pM3
96Bt3GmdP4rzmUWV8Jkyzk3Kwo16CDXO7p51qnHKZNGKZntCQJtd/MAAsjmT1XoHXNzDfsQ0zp2R
/aOdp+DMyigVZ3+YJEF2X2d6tDWIdR9ARU7zRZNDqLZ3Kr3iKTDM4XUp1v5vDgr7w9UEEBGH3MzC
N/08HBNkCTc4bwWVciX/eZEBg3+AEWlkuxQuQeDqe5L/uVq/CzsZPZSa88hZZi2/qd2oci1kfRFU
+Z+Ddw1SuTvk6h5V0+E+P9Odo2II5g0YjPaDsE8EO2MmOrajNYkA+AEjMNeTG3+3jvalhm0ITG/r
9NXDCNL2AkNm/ZHB56Tpxk9ywM4t4vrxEXcJV/v7WMD0fW5fTTTnr80//GdOPTIlwTP7r4IQWLqS
hjqXinq/1I/IEuUkYuqC3ak16hiFsCeJzQVylDk847r4NQqFmMSpj39bFdG2lkxw1PMB4m/Eajcd
I1rp5fA7cTmq3+odXSKs0TpWIeUUXvOA+N8X9kTOMFp7Nu1Ybb4juSIB3zrtN8WjuZ7K7bJIF7Ei
0vsMpto+lkCzjo5q9MaqGop/h7rcjYvpM6GZGHjCoAlL3vEUAIdtjeEDrFhRemRf958ToYLyPREn
3MU4+737Oc3aWKp2Ao8nqc3T5NAwtkEVo59Vze29wWmJ5MkMWQupamFquOGeEcrnn2AyQ1L6fMIT
cRhsO+D45lKt394tg6EKbLHVWGJH5RzFum8bIXV1s7miueJ/acn0whVAOKVq99jjVvjt+ZbJtUrk
6iUmnzeknnGu1cVhaPA6IMmPW8GteDwnLra2iCrwbqBWYwo32R5gKT4XKlxTbgu71VU+kh6B9bu5
iR/G3O2Ajwq+NKEMi2w8jMCMzdiyZq85GAIascgGzjpfqbmFu/QQMRyRzEaEwZNXkNKHRA0lg9Ju
CrbazPJtCm05wX0TqrBID5layOxbqGIhD/LHIq76GxAactmC/PV8Mnp6eVuWc08gk2GAqU6Cg5JW
mDiRJ770FddXgEcwmaGwxKliuCSNRZWxvdb5a74m/bcoX6aPUvruY5+nv6SaYzpVLS9xQ6qOrOnv
jVyKcg1Ipb7y4TuuhT9i4VVauIdJMacEn+KKzR1+X0bBnZJur4TBIS5AG7mYw0q4rE3vQSSKZoqY
B6Jy8yiVe+/H09e8BQ45XkplhlV4i8jpaCyjH5Zmeod0Sur/8XRzNbndGIYprwtNU/XJyeF7qF3N
TEwJy05+eHWZP5lMe1gdOcTmimMoqHs4IsMT7THAYJaz3GY+60Pwm9Bit5CE18LZ94lhaIXifY/B
y3IThpRZiza6bp1n9/TxXpqUqmFVZThd6jDQp75G8rLub1c6iCOn9Vb7jq+YE5euBVg9LsfxzgTh
uqzpMhn5OkQm8ZrxYp0AigoIuqACsQ+JzegV+RJRtp0ONHAqY6vqUBh4mvfGl1tD2Ja/Wwschf4z
pEMoycP6mouqrQGgFSAyo80zMYvrm3JyhIw9KCZoNNTMrwHnk8mzKNXSOSr6KAyVUL7EGazj+wOD
uJ5z3tdvzEjV5A72dLgoU5FwQ3l5Q2YI+xQZ8BK3OM9yyHQYWFiQPc5CXYWp5/lmODPgcvCD5aB7
GtPExmOaYZcTBOXog5UILzyK8426XvW9iTNd2+22j3jCeNaGXKrObjuzH0wQLuZQkjfwshIWiEAn
+R/ca1Kh8c/KB5axIwkbOMlV4oI8ekavP1d84LVSoop8fj9YXYekZ8MmX9H2yvRdeZ9+MdsTQQsd
VcY6I5gtVHjyz7JrBNFswvAa1Q4I+GM31zWS2Ykrt1Mpk8GpcpqX4eAvXlGF8uEx0CNu3Cd8c+pV
BRdGVVQBHisP/+4VRJyb/thThfhR41iEClwFZtoHnU1DHe//sT8FNwjqJ9aq0c+UGqfd/1/ccmCh
b6HbzgXj0wchmjQNoQOhREZY+NoJSal+CdEunBVWskaQIQd6ENMl+vu95WKEdQaBe8ELjhGt/50G
H03I/gixduTg3DDd71SLwpBg+J7TremNJAYlfpGM/4sn/5S1Fr0DgSLtgjUeGLNiPhEEulJj7Pkl
07qz81jGMFsTJX5BvOB51hfOkEOv/Cfietnlu4H31kHfIVuP21FSOUWhPgk++VqOyU0653xykTe1
M0zWDwJhOyXFhkmB2/h9MmaDmp6ZcsWuTx1vAYUgay2zRRwrgYo9XAxpxU5OG1XTfcDVf7gtxO0N
cFnj4Ta7ODxbD/iRTV2cp9v1gEcMnpvjSwJBZDZBIykdhnGNvXY9+zDLPp0RP19MR3ooE3zr1ls5
Yq0ShHJRYklsyu59mlcH7MB+upRCC9Oyn9tbxDA8uZ147ErZ0rWQdI5qodz13b8bUHpGn6WW5vpF
pGCiDdI9yk49QQga8TNTMg0N0cjYtbz28ButTtimbwb3kvFpS0R/2/qh5Ofy4XsKZjjd0t6bVhFT
HTjpZfDVGFrXiskTTSva2+aBNeb5npJ0cjwRxH7F9A2CnM0PnspWjBeMl9vJYdVEpY3YQsSNJ4zn
0sxrUZpk2w4T/Uw3GJoPjXcbk8h4hcps4c4DO2GOHYwJMKLECPb9+gxpI0UbvHFqmkKHHitLrXBx
zTjX+CoDo+Z2jieMr6sBmq+WamP0rd9UJGapcGpELIUKTjqS0r06hgzembJLHJKpODKEYz7f+t+o
e995XG0ZU8/oLDiXxQxp/6vQbhqQCr02LSd+nbzkTpWVnv7fmCqKujIPFriV4i62CwAphb5FcQc9
/miJX0pkgOnpVWyDTI2CCpApmuZtBpIXVaR1qfx4Ut3sc2Mw495iLFpvKfeixscMQDQhYdAs4z8l
Kbq2Ryb168BzoXuAA2ujcLQQqHnfQTTfeqaziaYpvIrd1OqJVKAIz9YMP0pA6EFX8BjJ27ijrhug
iHdeg2Q9M0bdCQBywRm06+0TCNGtKwtFGLkvitVdjCqrKyEd4H40t6Y411eNf7zmjmqeXzj7dFVc
9oJ6Y1ne07dTLUqkqtgh0LEtFDt31iOZ30Sp32TXhnt9OMOOSxbLjJKnlwP9Gq5WDXX4m7pwU6/G
KYmkzJ4eCvZD3ZkveWId86fpu70+pqx5nYBYsfR+yYaPCiNL4u/dz6FBLQKITfusH174ME63IwY0
t8XRuYzDIi4jjVu9z9bPP2oa3VxaR2VGCP7zzfbkv8RxsxnXgmXQFMT6eesBsxY54UVRTJwaUJb6
y/kIADeC7VTTTjsbvhl2IpNnbNty/vb0lCFpm7rbRJYLlTXFuqrGxq/1WY6eK2/tZAy8TzTw7kt5
gkQnr9WudSyVazym8y5tgbSx0rLqCHtOawAOSxa65DOKgrsd2sZj5cfz4EfBHQFvrc8DP+Rf8FJu
ZbSiqywML7qXg8J3YVDM5MA1E6w2BqtAsbtI36YRNV3+z0g39kUqnJ2ZPx6aAbruOeyvh8BDjB/3
UsFvf4/xVUvFTSfF1hAL2GIBFZEO1M1exi5dDOr5uXp9rqMHoLC24oG1P83Rn02DADo9FAbg9m5R
CcBtSza8rClYYxk3BvRT82ShZYRvXyzfSw9Srk29eBiJLr6+LNW+I0WvO70dWx3s6BJF+3E2QQ71
ifqYwNb5aS36+oyM2VNIakst1FWh62UUdEeOjNl7EABqjtDCB3dMjqXZ5rC39PzoU9YpzsRR/ZCd
5pmRQEBEzpLtO/te5FFOTqMahsgBdYNrjlO7iCyLVZviOXGsChHBLr/iW1dAsmIUGVJ6y7efU6RR
fdqQ94mGiu9HEpdSUBT5EIGSJ3HQPYs9EwGRw9rbdL2/pZ3FNyFlpAVAeoAwL0YUVcJPhFSkOCyk
Yay0ZGzjPb5UeYJl8SQwihaL7Lf0Ob3ePySXqFVcuBXraSXrn+afk8HU9KBmNVVvhhPX3gYtvvsO
48Zvxah2y9pgnEz3pmNFEJZC+WFahJua5szEQb7u2OQ827jJaRM9FYRnlep+CGFSUPztC18TJJqB
1lTilRTDiia0aXNnNFK3tpBePI/EPC7ZPqdtgRBOeGhrNluEg/taYAGFnwkm06AxS4Js54wP4hmn
j4dKA0122MODdQQez//50avLV+cXAGWYPilR7CCwI0nx5se/iJ6w+vbloXP5d8dCy4q5egt+diP9
jE0rnysZ06Vg+oYIOPP8+p716D23z8G24bnuEclI6TT68LkxieZ3QwErF272Nau7s+xw8ylSXS2T
QwmyCIYEBLWmmtbWfJgSUfeGEJnHDi0ZqsiehGnay2HefHkyMXcuGE897Z6Vocs2tOFpd4UaMdja
GvmapiY0gnW8ycm/RAsdEZcpf6dMNZtb3xUZ7WEYYu0Bx7xGN3nhbrC4edgbPAWGLxwxfqkM4qNi
+WP/gzH+mh/ckIRh+B8jytXCZXOTmTsjcmgOZd7Qd7EhTgVs6PHav5DVv5PHSLbNE+5YA5XzQN85
LKg0Bb0McIGYW5Vw4JKM0BPCY5c83J4en7j5aYIgtOyZSUBm5NzDWmSrqmCNvZygPfghN9vCLCYz
tbauMvTGUB21RMEhzu01NR8rSNDLM8bFaPQ/bHJh784rq/C+vuJMyMuw/9+4Ptte/FpRumOn3tGz
gm4qjObCqy77MzmmIUzjyDkwa4hYwBDIt5PpWt6+ZqVt7KcVJMTnwengvuKvCdBI4oEsqDmffdBL
5DyqXsEwJ53aFHW8ciGMMVHo+ls3EW7Ufz7lfq1Jj0iGrhRLjNaOrTgsiUZZNdAqSY2U7J6TSeLV
kcvmCpKiR/EZhu+toER53v1hvnvu1TV2z8jMAyCG41jkkufO0MLNJIDPE7Yvl6VuL8IjnnN2UDzX
Veb2rqHnlzzHW5J46hEqTMDjAmFvVcwOQyneWZ6VCKD0lX+yLKnFkcqBPyTbxSI4mrBO2ONNO0wy
DNq2CkswyuK84kK+nOMx7v3p5jN91PEiRrQo30e+cc4UmQzp/vlR9+OiamI18hFgIhYv0MpBwsp6
r9WGq2pfblJcYmLHrJ+u58OQhowqiUXmynT6FsJ7lIgiXskKfN5Sdron58/nRWy57+4UN6Tj139v
0kNpYMkk4qbojYIh6xka8VgKBQ65oIEN3aHQz7aJygHEGLG/nWClxdtKyqqlcWyIf+lLR1uk5SFK
KebnRsckpYH7YbH63rHQ7wZXZIWmo7v698FT+S6Yb7EM4e8YTmz4zpiErxocAja9OyCsBj/9Yq18
OmcZPu7jZkx++312CB0Vc4FBzwVoRldE9TAZ0NNBZoIaVLKv19jx4+kdsqusTkD6lnIsv0QkH4S0
hJjA86nGMkY/wNCnltUB2IER756yQeAhdcMmIRlV56SaT/+8AdGScw7wGJNSnhstqrY/9lurnrWJ
3Xit96tDtdaxndunlJBK1gvTX/urYTqPSFFBhrjx3cu/7KLUQvVmg7NhzRy/54wMLLL+UNoNsv8G
8dQuMYMrMcNswKuw+nOYcSkOlNnS89goDV5R90c4TMYKbQCwc5szvwNpv/VhgFJ3XnFOiszbANR/
WRQrIbCaHae3jXM2jBxeK0P2c2qkraEnrFbKClh89t1NXUkNiziXF1Y3QV5dfyRRdsNIbOGoJQfd
yvgWHo+qGjI9Saf3YTc8IVWMCYc2GQKbESrCC7tomyqNtjruP+MOBtkZSr8b/YHQQRQGuEEuWL2e
mDcf1DPkrfHI/R5E29a3NNDEWKt4q/sebFOPhCTNF7g8o+rbf1cE4+tno2ue0seNVfiC/LvOpsTe
0mi6QnKfpbktmST61hRnjLBrkdxYKzlBMaFGQrHOH7pS/rVj3HF703VXQYxWxupDDopi3vuPziYN
EN+l1Aahiqrra/dirJMxukCgmSYoZo4HHLVMLpRHD45Me4HYOetfW8oDTeYghskRGBWUMpv6vMoT
swvc7zTmosnYDxkOBCEPfcHBdAHO5FAEh2LpVhzLU6qCFcjcXLS5goUFycbNsG2L7mQjeA71jRFg
pNg0rvmdOIuG+JoH23VjOK14/8Vk79N9CeYsgOF1F3r3J5bwkdGs1CLR514Hc5QBCsaAp8J2S3hi
Rd/XyCqnbYbZAgL0D1O1JqGYp9nv/gDMBudWcp8zErkCiNdgUKYkATMt71a2V9SoP6INFVM4s0w0
CAuEM4H04nWNC8FTpkNRkCzzTflrYAjc5LCfPF3FUZ6ChFVJ596iHO/IUXd05rmvxtmX92APf5D6
dmpISVh/c2z10hHli07rIaLyzXCk+CwkI5cH9qT+HNPsXSOnO5Km4OalLekGondfX1XzJLr0fqw+
1zwG2ljNcWDPJggK344+nayRsaQlC6PRpHJM63hz5y7m9Ed+A9ukukuQI/JI9HllVkYydfwy7RPV
5a+hy9hWOy7+K8f5c9bpBp2vWcl1DooOuuVsXjbcsXHxKZSQjyOrJ0PTDbdOMXENY7+rWBps4BGp
fdYFu4ccUqgnTk1Ey5bQKR3kyQYPkPXq01cPg3LezXZadSrmwfUErpfDz1cItMi2ITxKwp+k5x7S
HpPn7u41QYCvaV1wtLCnd1wC18XAiJsjxaZddrDuUu/RHf1z+F6T3NnGXf5krdjo1Tepr8wKaXy5
W5YOYOFkanDVSl2twZKyfGGVucyiQ26S+o9gV/gOQH/lQNXj72S0WwcfEJjFmslC607RY5TN0Ddv
TBtEfXqc6o3xUaho2MC2aw5m2an39Q9mgBT2cdVLT0ZhzslxhX9UgIUd3rDUWx3fYHHm1enkHEQy
jtzqdMhbrXiXUdHr4uSseyDbSf0yJJ9WZeAy4R8jwvvf/8BDxtw2P74yOhrFbiT3hSdEUDdHc7z2
XVaPw08n5kB4A062tal/yz6RyaGEGQ6oF/Pk5uZ3uS2BS1MwPkXACS1+6FrbT/i+AdGqDqIPBm1c
B8IxOnIBkx0wVW9HzDGb2atVTUZ4j1uyC75jCKiboCwnTQhNgdenTUuW/X04IUIiGd6H5y98JXHV
3BspuZnDooCxx1ve/DKiCsq645802iWe/WogawHk+/gyiQoXrlCIGpKikG2n+W0i7po0TucT3NFa
MtSUodpHARgiumHEikK7UlciFaiOFc93UswMV0xueljgSG9GhTnyDHQuwKov0to2FFXVsMsB65Xe
ZVy5es2K6TXvJNJmf0KJdpXlwIhnehGbV60+VzoN9ZtWdkaCrJQLScVvVkJMjP6lCFrzPouaMhOt
MxUW3M9ndEexBEXNtCVLrBPOLmH15qaBVHU0bsuMi17x9/6w2GNxHde5JZEKNiSuOha7J39Vsh2e
z0iqtCisDSPlr+I9GM4Ejev+BjDWFGcgADAdmiIFP8htkV4It8JzaY8M9swIHUpWSzECtzOTl9zc
F+wbN/W9kdF1Z8HdpNdqRn6M9oWXP5adoZUoyLPGErA8+lA0+qMB3q8mJmOGj3m3XD6kw1k6ousA
Bme62ulBrSBPEk9uiIgZ5myp1vyIPigz6AkHDCwkt+BUUc2sRUBb60rdd0iFgNAdkjiz7Lomt1FW
XO1VdtKxGdQmdIDTjUNZ/AXa6RxhvkE8gJHwhgAhsqwHRcKyy14zYJT6zKqWEHSCHaPX9WnQz4Wi
CWnYIAYqOEroxxAWtOYJTMq5S+PehQ+1RfKZvDWb5YSgdInTYX55GFNbetweuaJRlB2vziONe98n
k8yldOLawHeAsTuMXX/lmdj8GVqmex2/KrFf8ZKliv0rp87drQrFZdbe+V+rBRHCEP6lptj4nNOg
b0l7cjCXRsUTG3cUVvNPSMgCJ3Lwyt7GPXL/emCHkGsUY0w3vNwRb+jxnaIqctMvFqRNVX4ciBmU
DcPtIQXIJU1ABBssT7yW6ucosx3KkIeOs2ZiZW9o0bHHF03+ri/6GkB/HbGs2ivZvGlhVI15Itg7
nODhM0jzniUND4Y2Ecuk5gRDuyfj5VMmL7z829rwH5kBItzpbGMPUgm3cYBGia2CowLN3JZHsvcC
vAE7Bxc0YtHDFbDFRg6hdRHfOlHrTdP16PLTqCM1afpSZylIA3l/QtqhA3LI6UqxRw9dEetdyrvZ
s6/gepktbvjNV67sY2EBkOf/AxEbTo9/rOXITIc/R6yqu3ThDqANR6EVd5PrM5wu26vR3qdJOuRG
ICYuECEAz3H1996xK61mP6qOYnoqm3bXThgfmiKsGFMPZZ2gL7w+5urPJxbkR8dHfklNF8RqXAdt
WugExgXwmjUXjTPIsa8nP8NkXOQKqUBV7YB5ttzDckvudZ/tqHzTm6Tr4Pki+izN5s1ocXmcSTjQ
qDmwp4scsQvTkIQQHFXk7TWuB+otCDWS9RQlAHFFJBQvHwn7AYmsoPbnWQ+p8y2Ysj6DcLzDMcEy
9KYPe9nc6+FUx7d9bdJauyw+oYgtOjJyHyfD6UBA3S8x0Cmb5aEoesW9529sHpJtlOeD2fycsqmS
hiBetKRlpCXw1kZBeukm+za/hPnsx1jdASBVJUpz5z+dydH00My9vJIxn7qX47phu3D+A27DY3XL
ocICjHSrZASxj2b9asnIHL3wrg5P8oL1WKEfN62teYtwkd4JboOgH1ul5tMZq3kVdv+UnkfA8q35
QCrzR+9Cw1+LVRzhzci6x8tuRUgIGvNrGs8ZjwfvdUbX6CzufmCIHXEJJgt24nCa9cOUJqZTCt9C
16uQWER2xhJR6FfyAXkpXzmBN8WQjrtRr00IjlA0Vii/nvsJWz655WRY3GnaoJ72dP3jsqIY9T2m
hNEAhFaVAuivlz367S6nsXwUwkO7vAXtYPq6heQZZzO3h1+s2KSqjHcc38/ek48RvKcE+DGNaVM/
G1iENfdpRdXnVNtiJxHJLgsPXagEU4rHGCRn8nH7bp9S0UWaySHNptUGp22jQaYSchkmXoT/q5YM
GLueCaQNYwk7qBPX5+qzbovWufS9TG4xsnCTISw9v/a941vWePcXCLdaQyCVVnTQylm1B4ZW8ici
wVKwv4sA/a6ai3kIlBuJdCZVamSI9VOnuJQYulBl0AuCHtPQUrYZRAVf4HIDB8Lb2iN2iWdbCigx
PqkWEpJRYVTVRMZVwk8PEkWzqQSk0R13B2hRR20flDtQM/7PXz1Sb17poXBxJGnlHHRFEBW1IZkl
siblH8U3nASxvtKysQrwJRaM9+xq/S4olKZoHRP/BQsPaSFE+dlgDhLfkBOcT9dEp7yKuoVLArOU
GKIN4NWWUtPvaUybIYrjUGrZNCtzHcH7bMz+/eQW9DzYuOYvmkww/PaVkfpuNT0IP2FSPmQ8/vK3
ZoxMD7vNxZ0e6/fjGUfwKOx3OCecJU6/CrMJY8HMaB/JPQI78M1+2pNNiH1A4JfsUzV6SXFfBKtx
N9a4dBFppyIjhmu+yqin2oGecEeP4QL04GlNcTtFUrMpjZWY0sYI2xFmE7iepuOGueNarKhKhisD
r6wNRskNcHEUwiqTCPknu7TuuS2R6lNk4xmGQGeeA1FYPL79KUyvGRyFI0FBKabKGv72zsMOAAG3
3SIzOfTIJbUfWvrwCQ/pOWWcXAg5ahAmpSyUDiWCn+3gHWlT7ZSnAo0tmmcz//2ddx+ZP/SoDC6Z
lTYtFGkojSnbbZBfD5zPU0zBmNlLrO1KvhW3NsLTG+4+LD7l8rqZYSUECXxpBhDEQa+gQb3hnPBu
Fu21o1rYxOa2/iZUbs0PAjjUHbIJLji0QWZP21fiuhjy5llWGINKGosX1w3nFNh7BVwBhWg7oPwd
Stj3lUTYnsHCNjMlpmEJ6D6YZ16Yxz24CabhccUzZnCAN907nvmMbez0AtPWH6cn9Jsd+csX6D4t
H6C5kD/11hsVgfm8RjFb8VgkUDG2eqksRCrIoT/y6+0ioQW2D4WBu7sKbmAaq8TtODNEvmM/0K/H
iAZPmszGjTsrQtq0QQXiXboWZdGcXtBbiX1r4NX6O9dhF06zwjm4TrPuDVJDWWpRh5w/2dHaLpR/
KvfPjCj9p70XU0srC1wrjS5FC+KjiveQznt+CeqhAlTQhFgK/uIsJpBnn48MnCAQgHw1+6WInUmd
45xfuxqTnZ3DrI9hMHF9+6wwS4nblChK2x3xom1GhoErdyIjK7cTjGhIYtQEr4fF+M6tiEz/mXkd
mzUklqXOYfd8JcPcvbutuywjMUdgQWZgJ5klvk5u3mHVsWAlsgQ0BLrV1ub5S9N133wZYoAZNIAZ
m+1xA1QHOZ8WZvs8Ua/HwP92D4Qj1L72LmdWIUEtoTnbMRHPRxt8r86QxWooe7D3OvqIfLdhVDLM
LcstXuFjRLxMfOP2ViUJJRrSpga4yS6Fq9L35Y/6/Zo3YvHkpjrZSJZujW07Hi20yWQBjx9r3Wuj
fDEoV6O15afwry5xJeIvb1kb45xZB703Vw0vQXcfR7c1f0XbfKZZn1osrgMSsWeo2BiV9Es3u/bE
+8SUFojCSVurYkdPc1aZ498hRd5ArKVkZY9cXp9H71g0yTLkOI6cGQkgcFvAP8MiBfjPlvJU9bdS
I+41/NSMFVQK1iWwmHe3LuIM1b4hy8g75px51kias3ZG8boB+rzajajGOh7zCU7UnOHqawEmmB95
KXBv0brj5EpH7afOPRuwrJcOrNTujozVwwBEOKhsW0PWoavNywrvfpnES3V4vC/5zBfzEoTCoqOM
oZmjzxgQ1sob7HQTl5M8DTWmvWK8nVyzMvki1TejSLXZuXk73O/DfTC6T9LUYN3lANK1/z+GC0rI
M30rMsQaVZXqrGIEkOERPJUswWU1nlwTjdZuV2fuJknbBp307U2OUogO4jBfoaub5l8xxOOwIeWs
ICI7yY7OwCMqXIzNUL8o4R0IRTaqsfVO940z6pekJmldIq0KPW7sRDadRIFejoXVrNyddyz9fo8U
D0GukXinpkVLoOVJMnWGCRdV2S/LtYwR5lEXpBBBsGO7dZQLWMO5gBzewE8SRZCaKZO6gFU/dtqa
gyUMqcGF7dlVsnrM6FKMuB0+M4Nc+qqpr8B3Yub4BEbwAlQOMtmwkpA9fNJDV+C8n4Bgvx9FQG7i
LTtttwniLYMTKxcYsTNrw4gTW6JZhSTcssJm4fbwNxWMNRdWd9JnsvEABmOyEGX2P1YlNTPkr1aq
NRHpOUiC9pzTDFrq3JhAcw7HlnyX7QEYbZBT22w1JB5PAm0+zeN2wyiDKmWg2oGp3de7G8YkEXPf
QL7v3+SdpIx2BhWi0Os9itDhiZ8MK2oADbUQy0wB4p1COCwHY8Nvdlhy677OeIp20UsOol/zPItY
2lG8Fo/BMCc4EE/F3fh2Suy3+ED4pFlTE8y9/fPfUUoh8wy+1PuW3LnQxDHuDlBd57ZkBLglD1rW
PPx3t/7cF8/RtjbTZzwBCcYLKBtfWP0HBPvlUp6gQ2b01Kb88zNP6xF9LYMTLdmBbvtBEoSDyl9n
fs8XKoPRLyZqHZLYc2W72sXZjhLjSjkGG/VYB4de4Wy4eAYd1UlR34f+tvbSjlHUnQISNgewSC84
2WUMXurY3sXVa05xtUiZYPhoGBoLCqmn2PEUT21R2vnB8i8P47O3I14VAbVbUbXjM9E91OGGrIfe
wgJOJ3EKP8mFjfLDnrQruUm8gwmhmRoAR8cjMZOMBjfnawd6Ct7+BMm0UxFzgzIbVHh4w/cmuEnc
wtePV1ZAWlAoYZIuaF3bCtQXlO+BnVnGZumS5XxIMDBoMchKKYj0cpgsUHKsnkkEOATrCw6rpLfm
YeWSVs+0BIWXvgYeXgTrBBeanAVVjfO67wdJpJ0Os2nHhNullsheLYxj8wwCzYt3HpKennVuPk39
j5PcLpA8bwLDqELjnv/KDkcljOD0bfnbey+TneA34Bi5Zz9DWaBOL+0xcHyoGnocEVGTUayu6muY
qtiPmM+yKOAYoNXXgqUKi8bKUYuMwXETriD2uYOplzJRlf6jCu95C2yPB7LkgpARs/zBbjmm8D4j
bam2IThBhPlkD+w5tjiUW5Gu13k2K577SPQ2oersVV22smvNOCboO5csozWayiodM2R1aM0eiTs0
6zpr5BrLOpKeM4af1cW8YcYfHO31NDbld/yrZSv70N4rRLHazS9DnKPqUzmsqjRDJJHIjcJCGDLb
LUF8f2VMEGAXrghLi4qnb8EsHSE5ibC0jDw1UzLcZNnsTTTzdrJJYUi4OCSu/7w5iaDCaLhgyPnq
cVhRiq1fk2MTvQn7cWtFJtHJQYuST1SgQh8JzIC3KDYndCRY3md4c/Y5tF+dTitrjdvgpwfrwYcc
u/Q2sXlxuY8rvup5RC/4GSIvK6RIAsBtyFia5zKoVJGVuH4jnMY1NtRzHErsPS+g5zMKDn1c0IeP
J4mXN3AYwd0eAuUKc9rvtcuwewcbCRfctjH/33flfFQ30tKwm5L8lZmKfV7PACD92tD2Q1pUs24D
8ZAOnVJauKYcRkVBer0fDQ1oDAxRy4K70cbGf1OhkObvHfc8CUOLVKlUKPn2pkqG2dphrmsT4Ju1
QJ/tCCx9r+kxs8Pax0lQDlLlsqk8fsEnbgiDOosRe8I5ivyIwLXlLk9ZIPlZoXLVS1Ug5Puxa+wC
3JWiChgwr79CH3gH+TGvcdoCJpGqBZbx5fa0gHg3VCRUBN5wVGF+uhtx3YqLzPw4oY/mnCqQf1Wm
iBR9yjktOjt6UR3Ik4XHOo1fb4zNJq9/JvBccQIpZ1DDiyCHRtC6eHYYuK+JcQQQWUl9PW9NGlaz
4qSJdbrM8OVB4PdWIjWQ9u8nm82p48ClVdr+NAneBQXeadh9tYcqBFgnlVzFisd0HhSn/NN/RE1L
wpb43mhQUkrknfniPzT73B9ZOT/j9jqTPwTtU+eAU4IZjYXq+CJYN2rZjbWUXlV1drOqJWyiRX4a
o7Tx44MBj3Y5nDJ5x7tCJcgiPVgap0sQ4DCvyYrIVNVHFTiutoWoR9iIS61AHedQajMFAdRVf7/L
KTS5xsskQ/51qCN6qFrAAWbpCeAhIWA9ISVrqwTTQv9v9codLaVqrCTwGZrszjGlOIoSFKpl7onM
xpZ+doadCLR258Ox35RkWRdKjGK0DBSXZyXzfX9V/ZA9XVlTjH5BKqJ6AzQRl1le9QuS1DeoAnRP
pvbWi2UNjwWDNQrMblwM7SmN03yXzV+Jd1ZimWw5cNA77YD65EPThVtNyRfVHb1xaPHZVAKZBPIl
AuVyEu8yRhQNme443v9Uu0GwmsjaB3fsoPh/fD25qTTkijS6aRbLAuCoJLMuBQE4jykcvZRxaCak
0nzQ9SB+vuxFPWNJ7uzRtl/QdzdBuEEnwH7j2aWGmsxSerzGYDsvQ1ISyjOhD4ddnYTit2/8+yQw
zeFgIlyyP6tTzE8TJkMm/lsrk19U3ckUJ1mLZcUhxAiXHg2xht5GLhAFCyGzr4jvTY3T9+zkPKaF
qxlMDsdI4acMERf13vGKhBKXoJZaL7vvMlTHjytzRDhRzi2vWLFGiRcWtyLUkPj2Wby50WlvdDxg
rbKnQ3kuVmvIAZYPZOVHA8rsOA+8ju9j0Fh81OGUqTJBpiIL4aEJEYJRzS/8D6W2lMr+KsYo+8uz
iaMfT0eiuFS7WeHVhTLQdBY/q6Me29G68fAF4+5wleqN38hUdd0UjJ8+p1SN1X+CKi3qVpCJ26O6
0qIPZYza5fVJLCmDBd/YYmjpH5nD+1fzfKy+tzpcZLBpeiDgH300RagMMgt/qmG/47POM1iJxf9C
EJkCoVafvI9oGD2+IkJ32h8p6CfGlqnkPgP9PBld+qC+99zo11mRH5BsKrYB0Utg8vcf8376o9XT
pWwaL+nZQNvKpGdO59lyqlbLJVwpaK6KGlIN04yB/Kxyy3nz1gf1TGA/eM6ps5rSreJrbg3qRvSR
cv4QkTh0iN28SD7gxV0dWHhTQpCw9e6WXsDWdh0+goaP4WrjtFgHOPmUanTpb7DgM4IOq7prfn7o
/WRGkPDbfwZp5RD8NndkMmKUsZax8XP6Lb9J1TLt2XepCZF1GEGX7/10yd75qdKd2RZHEDpDR8lF
kWskUXNHKjQoYHuFCwIfHzvmuCK+wOBWDgf1ywoGkhmT3YfbMbEX9LhCVmfLr3hF3eyIncX06aQa
WywTBI13o1jgIhkKo5b6UO7dN8f/GHwVUqwXxvgjOZxVMw3Npdei3RZ2su8VhLNT1K3Eea8nBqEI
ecMZqV7bW7U6hiq8ivzhvH0CxewOCOUZ8on7eKwACmVvT7eYkOgA/CESIbF1ChtXAgL8wV38+Ugq
nasl3GzmKl/PukwaBGLkSvaaKQa1AckKeqfU49LFtlwepXrI14yz6kuNZUhGgNmnpLRFubAnHCnv
tmCuOJIXHf3LYKG6JD5SDTxxYSbqLufJFXQ5V8fPQ8uxmgT/j23cv4JfIATn/0n+B4HZ29MEHATg
bUFsst9IB9bps4cft7SQLZuekvCUbkulhIdkORguesOX+Mw3uSaWbmN18BeQyVCmW+op8TTMmKC9
EGp562rIPaxFHCob5hlTvr8v1Kd6d2PCoCGtgDciDBI/5AJCytLQ/fQrbWnyiN9hbqteQ5k04Y9r
k48pHiCBxmB0AQA0roEzE+ppVzlwrLRzsC3LB7bxtkVMWu1u5RtvGXHyI13LOBPn3/zyZ/NtKnbS
lxC29qTtX1QNUfyA+RB6iHzyImpjDFiW5EuxQtYrvrIBK5B7fo7BTqFgjzULP08CUzLY/7m5WHI1
goeZySRGQ7CJk7RKgYzWfmIyIn5lb2CNnFhzVbyoyq8VkPaoiTAAwtLD3FRjDSfxyHh4VlglHnyi
J9ysm0o6990j4OSUzAAGZOw3aErwn/gQmF5c80H5mtoTbMZhYWb4N8bFUpWlZpr2BZVhFAyXXHnY
EXsxNxMZ3PofoxFwW68oukGXOtxHSmYTlPAxIePK78eqVAz2mFLWuVL3BBli8HSG+wpzw8sdysnK
yJW/RA181nszQAhBqACgblM9X4AqK9aBrj7oVSqhl6blwNyKe6tnH0BWDPR/CaPGzsfDb/o6gmlr
LSgO2XLqWUSUfnBO5XpC2Mu6oTBLv3ilFJUWGHruTEb93bIl5SOhfCDBFguhhLcyoM/CPUbp2+0+
2KqMbUNT7rfnaU41f7qSyYVx6iDzQVvhpufG0ycZObRJead2iCFKeuPuBvR0BnzhcGgJWxp3A+xD
Gs8SPA8dE4RSxaHt+5siuQsfHxSC/R+fbAlg5oGXHnuOk9zTe+VF3GxjzRG1na1Vn4bIZDiTsu1F
qVuZIfgl+Kvckra6KJe9qVYEEy2RFmFTvHLeR0vmMLCSB3rTFiyZyjsuKcF40o1BM9braohziHii
XrpdrvuIlUIAScKNA1r1zDe0rtO+2Hfex+lB7fiHVwdpT0C5Oypo6jUkfiS6/n2QHYUPSsb8eoUs
29HIY1lDAX92o/5E5whNDsBojYRAo0UP/+H5dIDGNND1Ne/5/6fHC5lnyXFzNNlo8I3mfNe/H5bt
xeetmJYqbNthWdDE/i9B7Nfn1HnUO2G1utN5NQrKYQoWcHD3QpKqXllNwB7WxGyZjLVbFgINFPMf
Q12l0ke9YZIklfnrAav8n3sv/RhJSzilGYuE4xzUXQ2B5tOp377ekG8Q6yP4mqFviMnCTlL2zgQW
HPWD9z1giihV29WlpBoS7j36ldheelJ9Un4CJWc7fXacDQcdNKg87Py6GIIKzct/mHM4pxbRgDu8
LZWN9fLMvMWzPE0USNrDRnY996JGQcsq4Q1liA7HRqjf+Kt+IXOpJkDMYMmbpbMRc/3xaifyR+dp
5X/UcssPEe2ZR7mi366zsmFITvk99jRJdQbLaU/Zx2G+tbW4s1MHDh+Yl5cC2hNViSwY5Rz8zilr
DQXQruLwK9fqaWowg9b9JbMsF2SNr9sri2IjR67avtHbSyleocs5uLFFnSlMkUfvQOcyjKV90mfL
vADUF8rFMIixMe+EUtcanfPZedkM03sYE/MhM0yGANKBEBwh2BxfLUrtGsb37jj4QuhldcRavSiX
ejPehlShoow3QTIYQl6sT2w5zCipnospQJplhEFVRIGcCa9KMQFKzZeNRO1aZVS/CDt5grU7V5hp
4U6l1z70qYhPEjwKrpXm77bt+XZjhGqfRJTB2ID7vukyXUfV8IVblzur5jBFIpEyvQt32LW1A5Q2
EDgt9P3r/3iaJxLF8Tl1UY5S1AcPUl3sI60LrxiDjEzXeutWWSGM5i3/7atvRJphWzNnosVkmVvK
Xy/bozhAnzIHvJfy0BcBkFSmS4gCbobek1XCduBI5y99fzLuxz6x5pryJl9Il98nWFNn10thAaio
38lBft5AuqiuVtNRRauN6YIQhhNBXFzCbh7OWfdn0jpqK8JjjTAvcu9eBlLBpHvGndHg6AyfwL50
OPKuu+OBGlenJvC++gg/dnI7WXnlz/mVE9Qj3PeVfRrbXT8Jm9uoBmZhCn4dpraBJRKkBfm03MKm
YJJyr1Vpzi0abZowVrZ3gv+j9Bc0+iIE9WtrSAJ/rESt3U1j4InEajFdxAcZq8PHPXiE93c4dQ3m
g5I8d8isNDPJn/FLaD3vpPpXBLCHZ33EgSJHK5HVEtDhhAPlTDnvJT5IrYPpoMPM6xOpo7HsIuCf
Z7IuJXctZcj0eSnMcBx5s3ftRVE1CAiTU2fd1ZJ/epRZCRXlzvzJfA6Voluz/VUH2nxM7FmGEA1C
RSmYo8JNf5dI2NiARpZc/v8rq3EcvNAkqSyuOT00g07aG3Rz6U9ZiBsohNGJswViAPkOdq4xQSjP
y01NyJDsO5KyNmFgJI/A7TRsokzmbrn5q6D0/kVePhaGbQaVsQdtsFiq7a6Oq4bXQj77TwJWD8Ez
im5P/DFmNhmQ7jHAHyOSDSjTPPHfbIdohn7d59MHqw0uSGmRWmEGQEJK5fa/iJ1gdoAdUPWirYPT
tqm8/zwPDTuMCrLWAOGujA/hpp9cScNk6wrud43gFNo8JPjq5ICkLQs4XpkNAbHH3AI9Sq+ju7PJ
bGZpCiURRtaJmrcpBDDuAyowT7mNwLTvfozb4qxsy215Weyee0mj5XemEyMPsGt1qDqVDQKCWAW5
WJH4BG86YCwsL0UY3gRJsX6HfwRG1ww4PUFi/eO7xclZOH/yoabDwUwnaRDCWQzb+03efe9H31MX
mZUNyiBJUcrrEoO04VIO/ODZZ+PqWcQ77ePdQZe+9wjZC1gEmFpyIpAbTgK/kKbwfNrhOgoWdg0D
dZRj4LW+JyD4DeOh5CZI2BkAjCH4/bU0aqytP4Dyarom7XTDYDdz+QTfzMQO5s/n+Ug0428BlTMU
cM1aP/j/A48vVwbsyI6amyk32hS1dOqDH7FYFA8ZS7D6xRyciYp7kJNWIqAHTlbYX91h5XqxRQGf
VEaVN4ErO3xY+xdniT/A6BWmMi9DitXFE5zilO0NOpTgx598AIae8XBP2jCdEBUUjmGHfoDb3c8t
PokCoSJviUxTkWX9t6JFo864McUGQnqIph6QZfM6mvA6G1/Vw/gcPjqNYoHCPGdKERTXLY4UpMlm
KT9A/wBIZ44bCGJc9kLy7m7W/haKhMQATkIh7EGxdXzm7fMUJlEcV5BvgLXiYLJ3UfjoKUmSstFA
2AETiLosZdRpqs0lApxvjtK9yyoJiLFQKcNBeRS6Z32HCDZIjH/BZkqYt964YjZ+0kht7cZL7cDn
cLsGntXubSyVNJ9uFnV3k7gGPPs+5P4Qc6L3nbsHOOiMTlPESdezAsfJFH6wY5Q+EBIv+ABnCcMr
jTDiio1UVr1fa1ipgJetDfhbYGRVoII7B23zH5YK/n/ABJQ5M73Y3ryyfu87KWyKBVk6Z5LCRSp8
4agfvczDdtpgHTUDG5gL2qo1aWgngNWb9ht8PdAmbUAdrIlEf8MVoQ/OLui3VEimpjDCdwGqol3h
J/UAA8MWoGY7Et9McAZq5U7t1S1FAIhuUsOi6GbiuBNwo/bomchWRH83cSMtyFotAY9PRKyRFsLH
J7bxHr9L+Gmo34LwOZAKyPxhlmOGq2Y5Rg7VATu0A1u+Q8w0EWuNzDl7kbaXix3VyzR6a8y/qoUN
WcMSB6vKxu/rHbstJwiI7j0FsoEFVp5+H43rJDH5OSgsBT3liemvT10PIJprKIeLdZfLMteJTalF
dD09z56MrBykrEk8X0O4c64vSsv2POwB0ccyifRQ+0FpJb0UYlWUqXv8kKTb2MbRYwHl33OOqdW5
wuOoknwh1gONeHoloGIvcULe6tqM2eWRFblbuptZwXxRV+MLDoOM9Dzx2oTTbD2AgkLIvpMGZ7bz
7zZkaOYOlRvuj2JAXjdOMU05VlhbKSwkIQ+AqBUxDxCtIhHLGdkNOLJ4Ql0qlDMP6OnmGrrpVcKd
CJMtHi65OC0izpNOv+oHGkCZvWB9Rd/4NAs6KbCstdobAdgowZANb3Pjv11tl3Z/VYKeyjnlzN9O
h/1O2z5vTy+7busoKbcGGC+M+EiyshEyGP6lGqN+SEuwiTU3iC5aVVPVydmi1N4pXY040kSpcene
0mplnPWAWxqeZN5F5xrrme1Uph5WovY32Z63wIS65c3o0Y7qpi3DFmrASAi56DefrR2OfAuBPANa
W6uVVUvaAni6tL29u7HFclqmykhTGz2IccT0loNvKq8wrclnDc8bMqyT463kzQ6rNfjiSKgowWyD
ycbnwnfyOhJdWxV0shhBp/1VEUetWK0IOLNHDUENlCpXrMEhYHQU/gF0vG8+neXwJanDnYsvx+cZ
X1fvxtYleHUYhAjmTOE7b7L8LZ3yf76G9p1UU8zCOcoaSB992vPqBTkMVBLkKwApH9/HfJ3rOE4c
imzdIRUigJqBrAWleeSZ2Tw39uITyxtEhPMbNHHDSUvRpNM9Dy0+31Xb5NPbK/RIUpJzIuDwbgKJ
r/ofbXylxMeQolyavWkVfekwaXKUP6iqPUNP6bEslPbi7g3bd4PeUyYNITGuO1crnHa7MFAXL0Be
4hGGsUOdWPutAvufO1eJv6fXHhJ7SE5I5bjh8VVSumSH62f66AMXtVAE8/sVS2hxNZYh3EfSCWf4
ELFUVj/UoUFRNSsC/AyOe9xhfDbtJeeb5yn2sTYYhz6cDZNQLFT9RK3Yzbwd1STddaNlQKD1FIl5
s4Nv+audyhUTKUdYEW2ncdh474ImzulJY7GEdTDg5kVhdSr74Hwn/ZKjpwtPBulimcL2aqZkUFUE
ul7r/dwbBWryY/XBhZLhYE2+uYjLab9cf5V59Daf0oMytw+hC5G9ndk/qbQvJzKoq8PYv7Xq2mao
HYNGw9k55B8bTBFuF7OUiaApAI3A+V9T9qq/UazwTCfXeLTPF0IWUxNxqQGpdQJxSbcBZSyeZ+8H
BuXBZCCSgl9DBKXfUUKqnXerPPOgE+v1G23C1HzZQoti37ieNe+ky2VWCZbwsKRRj02siBXjYNnD
UEtG2dewd1R38q4L6a2HXopAsDnCvtK4BqiPptI7uN1odOA+9yY7RnTTqsTei6LTk5TAUsEe8cyF
0tksJFGetGqv7Ty4wgXperMws5G8WIIMr53wNvSXIF1FTzWGd0YRx0jHdjX6dd0sFgFP9XSfdXrJ
gcDK1hjAFYeaNYFk5il1FEy3dr7nyg3lSI2fKia/czYnCiBfWx0NP8OHrErG1FwSkyiCtUPcOuh7
Jf6wKjTorVTkWNh0FGsNKvM3uNd32MHo+4EVgRQur7MmwGFV8qzmioDJQxJYxaUQJ1VVfqMTDozk
ezIgexrJWcGtLmvddSINL+02AOEFkYngyNco+moqYkDKBNB6dyWhVxwiOhwlcAB3t0pb7VfYrwFp
+BGq6Y5zQjD6c27ibgenFBVv+JbvfntBGfmV2LtWyawXoK2+sH0uh1jm3meQeX2+x6dpxbAQjDI5
saWfzqx2G08AF29O3gS+7lonLsocggc19fpXvyQGpvGOGtzWN+L7nZ3fljU5HfA6/yesSGPrntJw
AnZdUMpyk6TWNvCbx1SyKLSTWG1AERjyZE9pPokdSt7j/YWTvfCsi/yAnid25rhacqAcHpy2B+yZ
n0BSz28LaauoABwRBS3uCDF+fKLzlECNkyfZGAbjUtKCFoVGhj7RvQHxmzLrL7pBmxZa/z9cWbQ+
iynxNQstD9BU5wJY2bimZsX9c1H66WJNqD83Wn1itefVXFbK7S6j4YICjtOTC9EoeQQhMw8Ca1es
T9znTmP/ULeQthTycthrg19Ub9hIsG1ST80T65RI77jpi+XoEZdTAZjtzPspxJMblbDZFPNaq0FK
ySLxpGlUxryvFQvLMFtO4w2ZhGuDDALrPpzr8zy2jeVtYNY2M3LivVUUIPUNk5sv7g4ZYnSYSTEK
jk8tGVrN47aq0yoEEdZVBE1SFIAQlEMVmICnE55itE2cw/2FRgexDDUo7NEpxNJ15ySxAEjlUyBB
+d6li8QycX8S48nhl+lxBwf+zSNHshDRVYQaC1R/9/AaFcy1Mvh0iR8g2Rr/M4xPnxq7kcvAXp74
/tS9HFr74W8FLtJFk0mvwmWb8oIniPEXXnI7OqQOuqcRXbbKrpbX1K3/FgEVDlOseMmFSn/hS9qU
pnvaVAwwq5DldCvxWozuqPN5mr4zvuN77BM09BPhwi/RHaAq+ML0TNSkbrgmUoOkEYgQut4cQx1d
so0G+Nncwytr7wzsBP0ASy32cuMKVlDR1QpY52dB71z0ggM0y+tAzxB5MnSelyJTwvYeAzT1SbaY
YlG2d7hYg+5Y6CFXuPL+JkZIPEEJfUhqdArMjuc8Bk2cFIDfH0GKC2i984Ynuz4S88IAKkYLH37l
e5QDQJkmiAjbWTioIwOQIJlF96NMRsDDEK83y7kdmeJeaPmDnfizMI5m6wy00MzUQHwRHEbFR/g5
cpZA2eDgzPvzN9seQO0LI8tL2q2086I5qB6hxwj31fQOBOdw3yRn/crQEONr8gCcziqclW5Cruua
pqMXWKsqPz2SYDwtDsMWiyQVmMuDvPOrTEcQUFqlx8YiF99okuxXtFDC2EIW83v8CDOfNG6HICsS
v6lMiE54BkxAnxC1wl5VZVlCak8cM7S1BQ4Nigr3tLe8uBYX/T0eujlMEBZXfSpVsAs4Uw06r9Jk
+LAR3pmGpJI2b6Xh4oqWA6njBl4jFoBtLm+KQSMtWYtWpffOu1gJJy4guiOo1Kvs75JHFCl5Jc8P
Gex+2mRMe2kbKHmSkFiN8JIDiFcElL956jCa/hMyGr3YWM4AHrToAxb16l5jCE6jEOyqJGlMVWjo
HlSGESZZSY1T3Bpf9O7EJyLcO9+B67O6nHcXqviZkhbJOgsRtHV/GObl8W2YpM1KWUEvpPT/sVXo
3F+Udh+BJaFPxA1AFdWz39PSEwYUGjN86/Nq/6l3dlTeZcOwdqnl3AjlaP2PFmzh2EI28iHVU0N5
HHDW8K+9g6N9wICsJDN2Clrvt7ZZdI8hHnz2224ouLZFvl8oLQFxWMgyFZ57/8oV6xFEWHT+KPPH
4m5z+hEZg1Z/hzCmUUw7UOke8yI0gMJlAuVn6so/7esu0subve2XoDtvRHJpraSS1THbws+FmCvX
8eokmQTfSqreqSV08ZIdIvysyD2Tn4PpdSiu7VU2jyKmePKS+S477HUpCKyCtf8Ch66A2WqpKPfd
wBxE/7UMfpZ8SAtSoYZN9aPJIF5HAFTqM20HHoHS35E37FXVAstHEV938/1FHncm0jCQq7uAaN/x
0Q5WetRjLketDXL1OXH8EUDxt985ZIMEWcZ8SKP4HgvY4odJGKn2EmUNIQ3p+d1KyiZQyEyQXQ9B
8Iq90oVQBOvhJ7yOw6oILhEoM642lSnvFQS5324SfKLGr67dUnkJKSTsrIHeNQxntX8QqGq3HdO6
UyE9lRjkPuZIXFXNccZo+YpGc6OoKrEjyg4nGoQkYRTbtWbQTAkePPBrXDKvr/bJMe4d9o09wrDA
Za3/oMqCotevwXTh97ghfBkeXMo8383Gmf+EiIArhbXxRucX05xnvjWYX65aHujzCvjOu7DPxJiA
1o5+ID5wfBDohAy4bSciYfPy9RpI0Jdy50ZCOF3sq2WGKV3jh2NAgJf6Czu5bNLZeymxozFpYhaj
iX3f50MVsB0XFcKGUC1K/GrWllkqrnZ5+PvmM/Kii5JcZMPyaLVXV/UT0fBa/spQy4sZBQT+xPd2
iiYC8aoVYK2OKLK/8JPgPavoVXDbwXW7OuZya9igxW09N6nfR69bBLtFQTPmq1Q/UxZ5qAwxIRDD
cfeSkzdHk1rDsLI9COzUdqYSETfVXzJtHNMb/pT90tGdeHuYG11/yqK8pUc2lyKWHQCvryRpYYZa
iqztbvVIVt7sqUuam+WjVI7ZoZV9naSECUWY3+Cb9q3eBhHuvNmelak9vXiHlQt0gDC45MXh9Xjn
jazx6os1SpSLI2KHBzS/78iWP3aHGZ+14hVRP96NroCXTCPTKIzM1FP4dfh+UUPo3X/YS1zAhpSt
rdp3ThP7cshNV3/a2XaVA48rxidY2dZWXWlEOnm39oor6uBzURdQvjJMU6afObtPx3DkxyJu8qTa
l95X8m7JGPvK6q2NBf6McVEAL9I7ES6YWHTsOQbt+7pKDyGNEFd8klgKP9dhEKs9rVMsC74SNhMU
TKbu+b5oew8huHYbSL94hgx1QfX5+fOjCn9VZc5TD6vW7HmiGOfECFtj+r2tERaBIfkiHlT66YDK
e3wkH1UPvUVORdqUDTtzoiUjpX9hOyzcideYPUHzL1dARDXGVIiHsayuTuFdwElzpMiyXBqiGNEY
y7/Svz2PEgxLWO3TtzlLHDR7dJf2vmqHnSrHeMGTW40I4UKlvAThx7v2NPDo8Jmt7GAPwKMKQjN0
hv5glURif6c2vW3E1XOdG6c2K5mWWP4LM5bieUtpLWeHUdJGvR6XQOvak6XOGm5HQdA2e96enbqb
TB73UUMo2sMHZP7UwyUyieyk71UUCD8MZRXwKiEl93vq6SbcxlkqGGMWp2YZ9ceUFrvL3Ol86f4P
oR0vPJWh/JiIKvhiU0jt/R4XxeboSHEalTIx65FksMsR6nJl0XIc8nVbSWSiOvEbpWXyy5E3yO5B
6NC91+Nd/iE1Xa6r8O0F6ISp8ZuahNV0rwaKGddtYBXBK18QH4P+OryhI9NbfcJiSHxuK6HTPEC5
56+MVXUlSlTmY+w+KwTAJEImTA1zyXHxnJJUFEPMfTDxpr2cDEydlmvshXXO+7axzj6nkA1MTTIX
9BxBcv8jmv0Dq9Tja6wcDiPG0oM1q2YDdiYKQxpXRkAUdMG7sm2/Zq9UuNzXu8n3gvEW+CvhKcSu
lz+vH7DwzgetOQCwlIzjpO93g6h1K4UjbrGX8tLtWgaSKVk+xf7FroGB/jZcq++rkbS/IsNxehuJ
4L3G50myyWd4UGHUO9Hm+X7S7ma7KPCeahAXUd5EJRpuqFN6dP2dyF02oAnG+lojDgqE/9QAYcNx
tEAz7lKJ3/9TvuY89+iVWlISOL2npba0sR/g2Mcu14bgjwk99QpcsTYPo1pNZqmhqhVvub5oXxk2
TuD0d5gjDefuZ+eyiHk89GEqYNBJTbMY3EPEyCnMbSEz+ZjFG9EEltIKgiZyjwvoUS+s7IHrcOsw
7So7wR5fm6TRGPdOzm71Eenv4SDjYcohhXfcq4epC6EbZQbuJg4tPn/jlbH9WDgAlJA2St7gnC4T
+eYW/ng1kFgU59gmrSM3VgKONC9Bz3SQdazXQZeSelo1Qo+duSH/4ZJgZOnfb89pfzZqPDw8tYgA
Ihs8hj/DqtzSwn7Rcqn7lAIXJ3/anJlLN3OjSslGIVLosTOKUNy+JK8ASwBmSCmn13YQIMs+E6M6
Lflne0TyD9YMoO1gbzB06Lnh0EFX/NrSo3yUEu7EfuosayUKH4MPYupLqjjFUG0nJrj02MOHXMal
n65g+g8guxGLH59zac9YAD6NGb/tNexpSFRn8Fj0Rf/qOu9lIzs48FPVatcNrrZXEOazIAaJj2AS
4vUv+chs54mN93ibZVMbfn7STvL2ynbbIcYYpMGksoff6cn6z497J1w1DDKsMQiPn273Tdr17nRa
WBThhHc96WDfAMT98L0knnDCyBq5H/QYfrqGwQbhA9BPskqC9SjBjpQMJ9bb797PP0Lm110gSXHU
phYwIeA3TpA6oX/6HkJu1ff68vkZOO16P4jNHZkpkshx/B1//s124mKML1KY4Ydu26wiJy6Kmmey
WeGuAdw5uW46jVzcE/l1DQdrB2HWKqMdeFlAJdpzNXP6fw4L6lVWVfeVQOf9RtGi2t3EeSc/qGAo
c9jJ0oJTSXqebZjHLanwaTxkbOAf5g1q+oELsvP8hTYlnjB3p5qddx6tvL++sqNNxQWvfrKS9pVR
XUYK6ApWC6AxSIG4P6IbtySuPd1XQ0u1/iPcPQW1wDvl+jKUCAOEplPrdSesGnRF5XG+nJIKUE8Q
UeXOUAZcgEbNVD8tZ3iVuzdmxkkaZMQsl7TILqHNaGlmh8vZhZXP6bmYy9ha5K/wdynJSQ/5jtas
XnOnnj+WabdwWl4qFqyMfPKUx5P67BHE/GtJWZCoOlmpThTlMZKJ2OzkwtBmJslt3JmUXSWY4+C9
tK4i/BbiANmCbkpx9k3cHWyLOjXvt4g8MFAXeZY5CULTXmDwhpi0vlpdMoYd8+htH8tCNKeDXzop
ecZeGPttGRU9YW3svSBJRT02NdcVPA8mKxp/uDEcgiJdbuGM9GJykvKTfxVWI03sZ1h0mJhLb2Rn
YrxKPV9RvzRAYuBGVWJEcjk5Y6JKZPOVDOSya/37hl08+WkBhWULTympjnhcnwqLr2bLq7cseyQd
f9aGa/SX6vFtT+vKqRYeJ0NaDrOCQO3voKRiaRyNPgU/dsExQXN2dwpjxiW+rnYNjPMKquIJnBsE
VKs6MgnQHmlo81rdwDlU9cfulqUedRsfwL6n6gSNjTUdfThJmO6ZjKDx8WDnZzN2UylSNv4ZaMXW
Ic47T5ToQ1MnOoPJFWavOhNz/HCHJMdREiwnnohrRUsSMHWguGW2jsaJ4HbOELLdVl0rsDNlo2+N
8MWFmhQdbfeLWeEMy/FPyWrYvOtZK/RFLAWH2yOr+rzhR93u/XUoT4Bfhz/NChJMya30s5+acOkc
V/tpW2Y4m0zQiHt6T5YXOlyzWhhbNDahaI6l4tdJjNkhtXeoHo+8uTseP2Gp6d9VS3q/Ixao+vGl
DkMmfO7Y0B0s/rnUV0hHnycYefb4Oo5mWj5poLwKTMfk6P0HjTqp9ZFXRxl1qDIDwx0E1ZcC+tz/
8XHlvIXujGGwrodgAC9eCFtlPf2s0n90C5JM8ZXeZYDKXN69uAqPE6Ezh1j17uxKKwUQ5da0TrxS
o9y70+JMHPMuCgyAnSWiDfbFEYSsNJ+4Ld7oSxeAo7V64o6kxttCG9wMQaaEBJJ4khpr6XvNnf/k
EOY9sRtMEtIQZidGYxes5Hlg7ey2Y6Y6uEos7UiexFqOCCMfZPiYleh1ZKYyrA/nNP8rfcKfzIgI
xVimKn6m9GxOsfuvByYNCL+swLmFq1iuLfI1DgmeG2L9csWrfcc+Vlxnjx3iryNKmIqC83a4IcFf
m62mfQHDRyYKoe35u/6mUyhIuGPRIhTYjXuYuuCUPhEywDNNEfzsVMCN7XUwUvaYO3bQMrw/nfNb
JLDvy4LCtmSygIiMW6T5kOdU+BUUgv+C661fF+9IdKmv1HvYYO87S6HhNDVtAkItPeiNY7ZQd/bt
akjJGs6BcVuNxuHagtaTFhH735mHDyno0vaC5xbgZBIVKFd17ay5Z0fXjWuH9QnefrRqfXnkShDz
DpfgcfHyk6V+9OM6PYh8hMCgMNkaXKtuoCTi79kc1JaeE6Vn1STKjB43PV59HrhxBoCezZzj1yNb
114OuY2yD7t0fDGX51Q1NQpX1bozfICzEzP4728SaXFS1wMmUGn6lTovjVwubD7XQyuKvsWWAEkM
5Vt2r6J+Y9YWkAKDiXfRFS6CO8SI0iZbRQdGqbyKPxMvwNkxzku/nAbJAlFrQnranA3WaZocH0RM
FshiPf0d78W9rBSkv+PiJfLcSBu862purHmrvOyTqPKP/m1IBdnWuXXHwM1ALJ+08NdzokyJS9qj
ULPCEgGlEGus5UtJymGgHbbvy2Q+NY11N8Am9Rq8UiVer0Aa6RztpWKi2Diop0J1atE2C6UUlnTl
JL0FiWAO7y1Sa4vuT8dlUQbfIHq4r9mkOlSsc9i/fDS7+/QTtxOlIclJth01V3lbgZz/b9JfFtm8
TsUkgnrFApjJ6VkVMok3+2vQr3/uLSWZqX4nN+dCPZ9dQe9YUa7ZqhEDxZWOB9IosJNc6ckp80Xj
l3wL+qVbWdeZaswP2F9S2tIcr1jSD24s9tXjfX+TG55qyIrcG2GQS1YR9HlKB8b3rcOcix+IUZ5t
daIV+SFEO6RR0ER6fOkk+mC5pc2DvXGIUPQYlaxhc9vdS1Le8jlsOiFNHgzMTl0r4nAM+zRKA64u
nak+IBedCNjIyF8BkNCDG6cp4gdIQgnLhfv/fB4yRqHqtfNhGt9mt/opT2ziKrNC2fMPVRC/Ci8+
L2Ivxcw6Cs3w4ngAeoaZjmxD8BjBWT4LfDL0AMVH02iJTfF1nCQT1jHr8jyQqH4G7cRO/f/QdG6/
gUgmj4DYY1djaA++UHbVu/sXXlQ6czQ1ajAr+iGH/4zoudG+NoHrXD2NQ50WYZ4Di6TpcbWzKuS2
2HxIJ41i2DawAXpQpIuRCLfaGZs9CE99dfOttNlV0CXa04wdzcYJMBosSH3zFBaIyNp1ouXfK+eq
RBSheevgTy3xq8qko0UOjG/lcZWOSEFsBKen/ccVT0MgIa9rc9c6WxutVYdtD+h+V1TZMN9CpZGC
baYQgoEV6vP+wJgncJ2iEcuQQBFQmtUwnX8F50nOEeYHFP8bbhFM2lrlJFTaTZ/IuUCnQM9Ln6ei
/Al3SloiVTpv7rY7aqaVUnx/7KoS52gvZcCY2/JgKfpYqewpsz4B6Zj5xUlzBmx3cS34jb9wkXGw
RpiaVkqZzpjEs7xdkzbENlG/Hx7w6g9yoFWtpzKnRFTJ3BGxQFyxJyanJDplybglkXKkWfzjNGH/
CdHWj/7w+haysTaHLvTFF3+YznXgmzXGuHX1le38j2yE3nC7yzm8hRAZQ6Zw/cVRLTR89ca+Gw67
V191Y86SPCy3zmg3CzJ4v3WR4UfI9ra9AuzjQV9fZssxSRKiEgk2V+yjl2bnuqsko6MGmjPV0Jnh
4hebBKLOvOABUF/9w51HYx7KfdLZnkgWrpbbnGIrRx8ABQrRR/JFOOL9UVX39VvO2ygNzfuJE98y
gmD/DW/2xlPUikwWLN1EJ4dgvvzODKycLTArt6s9OQ7w44nuFhL1r3TJGtoElE24hc9jr434l4U8
JJ1gX1wIpJ0GgpAa6okt+QZAq6OdTCifPbiOTui8L4xOg8dg/EiZfUfdHYZXnwHPy3o+RbSdOIRT
FJ5eO9IrAmK8WLocIw0yD2ZllwI9jcNyKe6425ElgU4PEbyNmAriOOAJa+3KgBIodZC42zn6AS8p
YOVKmnYN9mrBr/yUbyQ/Tm9vfiKRMqrmQLqxPpLNQsX/3UspTO0iToO8NnQTgn74OG+Egr4sF0p4
MpAJGSoT0qwpTjCY7sFDOpFVqkEy0RY2JPQSBjJyESDtzFygvUqTcmK4iR4CpssIb5dlLHq6UvwB
vCE5nZL+eOBDjxwJeaWnxQ4bfv/5UEMk1Q76kyBnJUQVRVHcEPsru5rNYxGDdy9wHJ13o/aTnsle
7wLmiLUuooOvsjki5lWLPj18lN5E+WcxUI35JSf3BJskrNWtCuXLkvqs9hDS+C93oFZYTHGb7Zvq
X+8Swtyu2IG5l/EI2fTZJWKBSXvnXm+i69XGDl3Gzw2YOyeQYljUyziyWUc7xpzNJHh9Tk8glbju
wBqNMS5Jgk2f7dGKT88Dx2TwC28rESiD+c9+nm74TTgYJGHLwwCBDF7zhGlRUgkCHmrSVjPNkhN1
UtVqwjszrdl3PevL0dQK59Upqz2KfqBVXb+sC5uAylUkrI/OfXmE4ZsLOydYAs8ma0bkFCbkFKbn
Ytn0XZg5bS0hBffIKpFvyaoceiN34Wji8Nk+F5hdLPwVpi+aZdDrkLBKdArXEZioW4OEroLcB/aj
VYtUIkIJjNtq783BuI/envzjnC/B8L11dPqIMZtuw8eAbh1/CK0+TzyPDPMgAqR3la/74X6V0wpB
6ZvL7FQFlGhShrUuYIeJTQxh5vl8wDjjWNgDCnIz71ikUaxbXYODZmeYehOkiUHrYDxzkhePpsLq
6yeFoF/RwYcVwXd1AggAoZXnfetMIb4xUvNW8OFY7QLXXBISX4JUsOcv9nPiwgQU2wiX7FGwRNVU
MvAIncoN8Pa9CttOdOW0J2PPhLMCk4o4hCP3PNDD+94pu+IVXdt56TBrYeP7uqDo/XGqAHkX66HD
EKWzCprFGhgrZwXR7ZWhjv0DkP6/WpCpixtpd5ThuvNzUYXNalpZhtQMf+pRqg5aCHqE2Pkjxxta
TgARh8NwgIvEdqA/NFsUTlFB29JCzQlb6mFxalmRc9AY0+mgJunfSWI+MRN3fT5FqAfO8LWmAAaD
/OUhrhvTvWCWAolrNZG1c9/4ivcPR6WJHlbY3qVsgAYqH7yvwxmcbEwVeDIX4Vxyd+HPpDQPmkx/
bLV3ULyMaUXBagqfMcY/cz+Gq8w46LLs5o2GTUF9/mXJD5A3mFjYH8UK9QskPpIzJh3+ul3jTnFR
jFs5OzI4IQYpF3qBoi5eCxnonCdCQWJBuAiwENAuJiZjNvxyZaEH2d3m2+Iz5am4bAyybmPSHznY
bMyIJkxppKCqHLlxJW19wb8WAyCppLTBq5oFhPQl1cbJ7ClCprUMojbNAMeVJRtMmXR9Xeri4mey
RW7ZL46GQgI8nT49TAAGOQC+OgIi9a+87csNWePvTjM24+NY6MUR+Nh56iulgXMH9NQAFsBx5YkS
Xkp/IszQyhh2aMyjAWR2Ch7HVB6wlMvGo0zvxfFpiQqFzChT4dLYBhXsfUOBevrpZqmV+Y/Mrqls
gdinBZ32AG4azsucKGWeSlgKU90QnFHAgRuP5mBublRGLcvf8butGBZx1dKvQ26LQvghx1Mj8PfV
MrIE6+dNw8u+b1KNmK64IEk6iO3qphiqo1AohiQm6IdkxDqjqfLV3Z1NVA0gL94MNCugmG8CnY82
7Q1tGCYc5WXt3v9sVnym0XErV+zU+Uyaq2Z96kyjC5GHFcqEMk0DKAzHdi5yz8DtT3Zrm6T9T20x
mQT36lY5Ke7NAswIQeuYXXuRRW8AzT+Wrp44f3BgkbOJu8ZnGOGRXl7q2uaMSrQfo1R11fkeQfFf
sTNQhtUzyahZck4QFq6jXKNF22g+JKU8+Q4If7twrr7aAidqMc3NDxC3xr+G925nMQqWueySq4RV
6xbU78k/bIV7d6Yj7ODm+5lnjzRxQe4kZrPyoTE9BsNPJKTcgj03fFNgIWBprs7HgygBJfs8mAZI
0hpiYI4PB7kj4NI7HOvGpkJkwSxla65Q0UCNsN04XnbLNSjelD/QFSSqA4rKjpblzxSVtGPfofQk
8hrSEA2zQbT4jfFGaCDH9PaK6qmElngN1IfutjJY/NMQhaXC7VjPPbYF4PwlcDthNQdfoLLTfGq/
8MXQZJh4IBB3Y7d6Gl0lK3not6EHhmPlq+nJaNHLIddv2qplt7Yxg+P39ggK8fKhKh9FurLxbYK3
4dDUwqKj/w6JA/dDwPL3ZWbE8Dq/bmHnRi7zYBRE+qma3EiA0+cEdBIAqV/6oJAfDvWGCxRLfHPZ
3r8qL7wpj9nzFNp+MGSwrdMuw2IaTZAahaZ0PehYjNUYwFHVaIUb1Wz7pd+eL5qYZAo1wztPKiDT
BJS62Pd9YdGoaUfZF1+d0yyK1Q6CpK0V8uDCCgBS7Z6Kohs6gseyfyJ3YMC0Kd4sBKXjxBgCuwxp
lGLpgwKfpT9y95ofRV1NYb+I34fti9cUNy5q7oHewL0neYLr1K8Z1LUXHjNSV2Cb8X4mP/e8em+N
CPJzsqFW2zluTYc53tbS3sf66I1UUEE9ZJGAIPlNm8PM+g9pgS2vL8e1zOq8g00Rs48pVl2XwVEC
YbWYas26U347a23EM7y84+eYthAzbB03qO/aLH6udYvDQcoeOFFy1MtTG5sOg0JbzwoyC46G/TRH
F9RfxjTvkgn1jL63OJDRJ7KxH9zkjfiPIMTVKQFQvasX8DdMBcOXEFpo3/Ldu2AR8RY1QYVJmVbF
glbR6Z8xMQ7j14q19BDWDgsJNm/qyr954kkvyeDyj7EiabLiMv3vZ7iLUjgGSwUXS9Jnfzd8hMhT
6wkxVgnT2NDsq5Cb+86UhNueruY213RWcuyDKpzgubBrEO8BtTWpG3MmDbeS0E7O+jjZp66gNFgD
hblsms7MNpAzLD/dm3osIt3fCArln5RDtWoEltIuMLvb1QzFqWnYFlQ8rk0pCwI4VrcrLbGwuUz6
f+PAGxWxsHNQ/7Mi9il3dYloyklHwUKrartvM9Pb4zpIDX7XGTrGSjZkzNM9gbKJIv4SkgpKmfKd
f4/WlWa7qFptV1C5eb6KK6M303gvGsnwCCtkgaANnP2WVyy011po2AVsBtNPt10ZFxKOns8XU4G9
RlTNCfqGKfveSKwfKfB6DFz3mh1rEE6lmE2Za+2g/bO5p5ucnWkA2VNhceKm1QX8cF7nu1UOggQ7
bwcRaqAtv7lrbMtakO4bjQkL24xORTcg1YNs2aPFOpjqASo6IvktK/qEcxfM/YhGvldIJNsaJZgo
G6WYgcgnOEe5KohU88OeW2abAse3KhluCf3pvNE/4wLznxcnc4UqY4GCXzDK8MH+fWGffjsIJGAv
gKg/XQURXHRsoYNtt1COevHjLtD6FUZ8CaMJho0fW2Rmwoa0oQzm/b6KZLV2wBaT2D/FA9XUjV+D
7dgZNaVRk81wJQkl+O3BN8H7nztkNm4EFDWzjMhyY7RujFwCrM7WcczJhvzcT7ynWFqK536mfx9E
08BmJDtb6G0nPzv69VttOdO+bJsH2hVgwr3fDkdwWzCb17eh9iepr9nQw6aP3QfoUhNUf4Cr7HZz
d7qbznD+zFC0VZSPdQzOpvn8fD4eDFpf2mvT4y+Qzo3OXyi0iCLNTrjZfP7qCvOHHVxhGGI79dIb
MzZ/p98JCszf3agx6Ln1WclRAvRzh7L6XWCHt/N9+dsrNZs8daD4KpVqwMvE8MhuN6CBnxKytl7y
7mPpc1L2d0PjsXm3cEkbr+bwJNmInT27/yCboGzJRG4DJCstE4D7xLl8jCeigusPLOvOeYUWJDNq
VWytmaeY9ev5EkATtfQSigRHKs0TfeDQsJme1GxDn6n/2xng+V4OKJkQvPY9gbsv1R3YYu5YTT+e
1i68OxBLCjc+zhlvs9XJ5cZ9/hdIyc7QyzglEr3ZDOnC3iiEogbLVeiSdAURm2Mvg/a9gz1yiCCN
Ps1UccQOgDO97WOpiK/txKLSmCFMVvn0eHpvdvSx7FV3XOFWhs8LrFIhBcqDGqyWXav73qr2cGDa
wyT99XJmNE7bswwJwA+FU7xcDhsv54JAY8M508XHc+HO52K90OFeNkfzSFWxv94QGOE6tLg5UzIW
HRi2Wr+Rcnd+GL51SHOWFQvORtRwxjYMtXyJoHch0iazNMT1OJ4QwLtKZ44v/Sb2R8fJJO6wooZ7
GHFVmu1aLXndbr84JoVeb/wbUkjboMjb7JhNgqFwP6Qk/jQnGvB5oVguKuBwRkplZpdXfUBlcTlg
O9RHC68fkALQru78rv1HtijJMkw0gcWklhve4fe63Xem+z/2IvJq0ghP27c2PWvke7XRCW8F4MmY
NNFZGBw80y0Xsh07AaAZPUV24Rt5eHtT/U5nBx+rv69FpEukXearjNSv1c86Opgs9u9xlZYNotgM
fuZEKN0tHhyrCXh3qnkTJIOW/kt5ie21zT4Tn1wZ5Z5XEwCJ0OlPHJrBkTZUaxsEggaqDNyMDt4w
T76EVilw3RcL/q2cadf6TRglQENZD/DoYQ0TZuUhl/TyXzP5eWFArCiSY6ERYaCfS+7SkPxqOLAH
N8eTFpSWLJNbvavR0/iIplPmavyu8+2yOZyQNk/xZnvMm7oeHgqIRf2g0BKoOpfc6kU5Wdk6d7gM
4DRyKnW2EiSCl/8n5VdMdiNqEelC0uwYbSKeML79Tr5pquGSJtl+XWjF3Mz57SLP+NghkdGarHTz
uGNQGIwM7/QkhzT4kUrgC9oHLu9fvzhaacy/kgil1NWAMl84FUsYJfaA4thQo/J8GbOjsrlYIWNq
BrwHtZIioNo7OyYCAMa9kxf0v0TA+00WY9DLlmVUqjgLLzfvjXR7JxO2/aIkyK/2XxjqjuC5aFQj
MHhUy5IFyoRgx3DuAqm0f4xFlHCTNYpQQjY9I18OtdCp13bn0duvDFCxHImNfm8qVFCKToy2UgLJ
r4xavE6CrQ/31KTT7BmWQZMemGstreKhL5gom9mdE+GExPVkftIHvj+GpArAyDWdqKHar3PPzvBD
cNblJnvi1SsiQ2xuj+1cjoTx9vj3pBK7c4lVgZtwvl3Cp5udPcl4vtYfCQt89ecD008AwmyiE9Ny
OiFXoDkx5WRwA1uSWMkPi0LmJ4XK2JWNm4a2tbftgfVqyUaQ0p7XFz5Kx2lDZCWXcu8tEF9p1X4t
IcDxcNuDP4h8uXErvX1YX7sTo11sndWxZd7g/3sQHuyQ6/cRPuFQy5907fdUXrmVnysew3VcrAjv
l6eq8QKDNpYVA8cvn2bkzZE/2/QxPyVK7MMVUXpyDhuWpINVsSAD1MmD3rxmMV6mEYNBRUZKG16m
148ljOmNqy//at/JQLwdKwEOrA6OP6NwQPQ0tAK0isWCjh9cYUH+qvXh1Yjs7fJV+sncf03o3OV6
nLmEXdZ7fYCThZ2Mw8nC7UA5LoRFUJI+4K78SRVZrc4+UV0iqHxaCx5uxTicj9z4fsmZLwXWvj0Q
F825SRASmzSvMK6ObLJzL9RV3S9n9lhWjDMTH1xynjYSefL9BclKTpwdTMnxkUW88RN2n+kou2aM
t8AYd0XttTtiq4ygxgacMLwBt3yAyN16Sz1UbCIcSvxvamS96V7rTRFFv/Y08zTotNT4Vuh+iMLW
ICYGJ8GU5RJrONlS2Gal/7TY/4ZVMyxzDrrQb93nzHtbIGRHyFC2NJ6z1aGwlj7bwqQpIbuTa98h
8s+/Ww+fh2n+4NO7bqL4aUkLb1MZ2YggmxRFdb40x0h69FfQPOPYntYwgTeNbd3VG26tMz1ymoq2
igfgyXpvSIfMV/5PdEmmJ4vdozXBkltiDa2B83K2kv7Xls44qmFigkzkUrNYHQwN6L94K284jhaq
CcSzt9w9mes3iWzEH+2JXw93yB28wfjw2hAO74X8AOWJpuxhCO7QKkiT6pYyq65S+5HdgxjC9hMd
de8xM0eiY6pFvta9EM5LPDC6Ta54IdksDEMiQkwFWpP2aaEHtVyYitd6JqjR302PFGNDuj2Gv140
WVFt9pbioSmLGIjRI5rPq7mIucEfjhSatCMqnEtlP63WbpQiTHKBw9jyPzeNTAI1Ex+aYlmymEe6
4fhfF8yd7UUOjLk4y6v3mKp+n8iRlWDbpVLco0jGoXX5e7FdN1oRLRDfP9u/y2aUUHRlhkEOj6XD
dyH6FXq9HxZgvhhSwfrRLKcYxkVrH9KaLj1ZyXmIK4tl3RFGRG7ul4zi4itZ7fa8qXkDZfadena1
+05pibTXvI7UlikW6+qVwgbNqBFcJ3Z05UDTUf68fdjJDf07KxvBEHldp9mteS9J6jv43hxs6w0f
FV3xJCOuanXNAMEbtrg4a1MEyK7zbklHvPMLs8JybUyLJ2zks+9S0t8u0UkvFp6GzLW72I1URkeq
bGkI2/aZZPcB3XsjluQrztx3lQhYDOpCuVY0y+2NU9er7QYwwrUU62uTNjltEq4PBrJNXBwy6WRo
XJzqYo9PcZtp02ulCwqlWklsJGhHgjeb0Y0OB96eBrUVT8hjgYhf7cBEBb4D/9JhTkCAtfiZdAgL
W3l3YJrPIV2dTr2Qe/bP5zogPqsSt3dOXVO3BK1OGVtsM9R3+9HpmAoMAiKS/c5K+NDT0AhvjT8D
5wf3cRTsyRn3FCCrmwBq2kX6ocmWJfUFVv9hncJ/m8tOI+275ssC8y+jYT4glQdGeR/k0DIRQUxZ
VJMP3cD8mVVev/2s3hQWfPWeGrKolccLGRuT6B4Evl2ddkV59ypopoJjLPteSsx/f8Jrjr1k+jdV
W0jRZutSvmIiRPLFFHaU7eN8YjmXtIhZ22yXuEGT+BqFGX1m806kXEmGOanTZBtbHwiGIM+ruAi9
N6+iGnxN7Htw7lNudU3aIDAd59tJb/xqyeCrZF/e2x/s9Dij/njh2rICHTBrzPCgIZUsCLDMxC9L
71gqrx/dIAHwuTZ1SJQ2KjoHaqwBxzQrRGuEv9srb2ZFOprgFrDGX+dn1SjRxlGRw9R8UmQIiXY4
zMybqdcnCKUvWb1yo2G6hVU05UL/sFFzYmJRIARItq5pzXQxZDqal4H2abyV1cND0pwHlCbfJ0/f
E/XLsv+hvvnhhNot7FFt10eV8mkmpRK9VQpYSUDiwtFY6RxYbM9xuLh7/MMhI+ge1MUaX6sHAco1
iFNe3AoontyOZesBWB8zrjintyYK2g81AnErf290TZ8jgcVilV1FzJEDaUp+XV+DZVfIpnHYtxsE
9AHaEN13F15Vu0YgIA+WQw5JCydEUo36YjJPAuKVBF1qUMGFUkvdFVeKFiOfFdbGnlUvhjtkbclz
+d6UNPZ+AUlwewypWP1wT6ETKWYgSd6e3TIi7vAktOdKftjN86w0r4jaTxCh/lqJosVJSZuxe7JK
hDtBZgcwK6XGQJFyLvxOwCsBXv22qmML4AIyHmCLaZfK/4NQwB1v5Qj+BOyX9QdD7kFscF+EKrDt
MI6UHphCKk80Ttv5efeMuE0bP82csGdCrfe7y9iBnoJ36pqXuSu9cwI/tq7TNeB+YuPMPPuVBm7V
NslKRdrP8AfBJQFzKc0LhYbrILd36Ycw7TyeezHlXmf5mQF2LR4f9FupcDVwcgKpWJdeOh/DvSlN
Tiul6fA4XfMJBhSVKiDCUqiZAiYkqJtOWVkJNpNBRZ3UrWscGszVYPT/Wj0bjYF4A03X/7RqvDsQ
k2bbtwqLicoLuKeGkx3BeF9uaY2axohDmHyQ7gEsB6AuDdy4L2qjoy9Q8eHIe52LJnN9hVQIwFHn
kbeo7EpSW9or4ATIgbQUNbByfVOjykTcsD0G3dzUvCklYFMq+Avt13VaeM0YdYYHyBMmJIyFJ6V7
ReR3d3yJvbHcxaqeQThvK2N+B5QnORh40lKNu1ajGbaICHGOlW9CkzUPPSxUUyOrrtIyy9t21f+f
AmtsvIue277/PMbtPgtSd0CrtukR1mT20hB7lZcQvXotzggWGFsPm4TsZ8pPBWTTzRzGPBL/K7v3
Nvbzf8QvMk9QSF2H9MnC62/J707BqGbsFdqZ7XmdFYmOpAZIL2k4e326V3O4j6SSCix1EHZ7HHcj
oK7i2e43SjvbU/DxDxfDurAdh/pS3wqGg8Mg+wlI7TWQsjfRyyX2Aas+wi5N+n6nGcGGrGgt1Zln
wKLpMoMIxNBavGAckjji4b/aLYkyfc51bAJGflSVPQ8G4EtOOoOZpOkQpTvRL7x8TlKhm2LS3ILx
16BODNtlqF42KSgU7YzA6jeQSPw0mGSftIiiGkcQ8w5Fs3nR8sTV4lGo7p5RVTvkw7SZMi0jZy1m
qzyMdCCak5V5x5Wczem2RD5tIeh28iqafpYrmZc/bf3Gpkx0xU+VaeuR1g0wn19tgk5r+DCKnTXU
IU8Qa5bh1CHdVjixDd8DRcTCb2C5UBybRqTRAm1Ze8HYAhg5fz/ybOMTVDFmfetManOHYbVRdXl3
V6CbCAZf36gul8ThiHWIA4x57X1ISjTe/tv8AHr/WCV9B+/v/3o3LQLwXlw2MfX46hVPVfgX+bIb
Va9O8ZKqB7tpMCQlDoTCXB2UAxUN35r6UABaJzqYPl4IVxSVZmIMNAy0fa/DV5K9xsn96iQyB36q
mW8TMYl2I/eWeraS5LOtToJuh/yvl3IYuGK05xd9UZHy0+WGPyb7hn3n35uhFGX6BBoTUm4hTLv7
zF066fYkxSM+487tO/9M8YBS3ulkN1qzoT7H14sgPv6Jw2aJzPSSpKI0E2I/5e3wXSG5h1VYQzgj
VOA+YZVdngi4U9KfkXXMSUhph+djol0hSoJoXG6TeoF5UR5mM5DJwXSG7gaDE2LSjSJc2Nw7mSfh
zftQZ/haJifSYB5vl+jXuWA+x/m5R9o+DA6faIcg97A1/81Ehs67XEKAfj0+Y2UUV4gSnS51hPm1
UZzoU2VKEG786yyRNnMpzdUFgbdaHiXTDAteacvkI3u/v9Wj558koJaZaA5cszPw8kjUWuSERu1d
EJ6LH7v6oeuBYnTlwbw2snoyvSMy3uGLvVMJDSRsPzvxKmWMHsL69GgChgog/6zEYU/yBMN1JpYq
G46SQhpuH1JMsjxDi/NV6j9VD4BzOJh/KIDO1h8kTS1WOMBnmAV0bew41xRVjj3Z/dZljMyVa8Rz
lKnkCnaLeUXHYFOVScY0c+yL/m1eFr5Ri27vr9b4I9zRDfB4/hMxjz2UZTUQOXitD0tCqCmQLAEM
bdxl/OAUtqVoz6dWiX1jW+PFekT2PFQmsAm9iFPZg2ueqxYu7BX+BjPLEJ2ABGHnB2ntCrfdcuA7
8gKtxrVARkRIjUEzRqBrjha5j5KJIX78D7Qihv0bd4Yg3BF5Q7Aol4WvPfSf7ke62u1Q/qZxN+TR
fVEwmnTMzhRPlKWa/gP0U1J+fOB02gujikvvGhMnb2RC6BVTVrSnBjKE90mfpQ0OpdRCry8oshwc
xqxF1eN/irVeZMjkUAXtau7NrWDEYLEaOUOjMHpy2SNBfdxKSU4qrCEHYF03rpwfQx79uE+FNO3Q
deSylGCWxzI479qvq32c1y1qAJGFJmNdf+uFdqnmlYHZ3d53OgWXFU/tIVp2fT2iRiHzQHTL5Il6
fFvRRKTH9httwDTknomBnsP54N/uH7KA3yd2iVumjy+DT1dMdXz+bSjaFa6TBg50SYBNymhDEl8z
1ko4Z6NtsDW0uY2thH2TUOE8CboKtIoIEIzurcJYzmx8BQ0EW16jIJiLmHGiHHIoZCyDDEq9Noa8
sfMnts5sEMyXR3b8pEL0YL/NWVGh27V4VavrUVlOLcuodVFXTqVRaZPkoIUmnTUsqxUpLELBmgEH
7Wx4V0SIZy5hRjoA2GIeZo8b630zMRm9WTIzXmnMYEgV4Brkgyx+tK7tn+43RRyEcR00nfCXKRCN
xR/3O1CNiSxyASfPNs14o8/R8fBniA+XcMQnR6nhvvAMMAMLmkDuEcG1vEzF2YP8fOExNAMSa+0h
KqmaMUSAodyWHPxrGSD5XJXtVIjpDsai7Wo80vprGdj+N5W+zJYCfXdHK+jvojfw/X+3W9hY2dIK
qTFROn44W2QS2SGVI9zzbdtocHokM5xTf6HcRj6ZDF2CdQgSof3NMD0GHhzI5WMyUGxNEnUtZRFV
ybnEbTVeO3k9I6X64HWrjiJblPST0ur7w1P2gKa1Vk0HFTl7cEAKjAE4/VCDe8KkxcNdWUlAIyON
BpRPQIx2WfhtI+7O9EGzfjbcHrUOTiMY6iel3vatBDIG/NR1Q2ZzlWt6J5SEWT8DcZHvnin+gmyl
k6e75JeXmetKzxY74f7Y3j13jdrTiz/EJhpzFIgpBlPVKSYWY53PPvg5Ps5PN2NLxfWc5JtMIQEl
HkIWIJoO7EdY+qiCH+pdLZGqfAh85ssbgP7tCJfrQq1QqohyYHthG8iSGstZAGxEhwLB71U0e5mI
04cHq926QH/O/bePhEGWm8JYFbn4qRxgqXoX33Jtk5iEhzDSe7hn/AdmafCMPbJyRhp+rpzCuMvw
y0B16+jbu/MdWQ2Cd1Wh090vhxrrI7RaAYck1rdvZhvvvbthXz8L3vJNb6oY+WUyto1H8WjGcjYL
H+pV91FTZMVBsfKQRu5Q8VUuke0qawnp3XD1u3XRfug5JpbROhVYrJhTY91FrbzDbNZa9I5M7kYs
J1iHsQmqe8EwksTdSa1oVo3sVCc0aaHTUqk7Mkmkd706pHRhC0bXX7ZuXIZdzqMbKWsDhJzg0Mon
j01+8FLc3SjKosbzKCqKuOCxHp5U/oT1vsJ6EbX1b8ofWIQIIL6UhLaQRntJagv7rGqCUk+BRX44
I4xSPzzAxkkuzIv9T57wJ/xtcEhxO/XJAiqD2qC3iMh6DZY574aR8ygDjmA7P/JEuqucH8+2HeXv
O5UCOSUrF6Qlm2hSDp2pMqQ3pf5J08lnXSf5XSpQacGsmI/zHAaRl0Aw7RcNP5oPd4wg4H17LKuN
T1c0P0ZdaxXCjIqPiXLgPk9jvii8h5Bky4yvsas7rYEZsnF6XEGwX794zGefsw7LgTCWokIasDU3
pYvutKJGOpBgaRYeg7SectZ2FJYvQ0KeurI/y0YtOdp6/Y4wapaWyYgy2hzoPNyYngOpa89r4ONy
Jl6j7onC9Im91DAoXKlE+XFOhoCvlmeaghgmTwgkdxnVLw4IjAE0IarZyQ77xDtPCvsQTCv35Yua
QiHipoE0gRovw8IgY2nY0XWnE7WkbQFTWS6LSdCU54m8ydsRCFrgpmiPRrZbpvy/KJoax53mn9kg
oMXPVExONt0jwZpOpCawZEqFW1VF+63HLMfQ7ih+7nEbePQk6ZJgWQX3bn/fVm87UZ7YkfzhdkjK
fUWAGJ2ApaM1W+WbeBB+l8z6rj85n+HqTzCo0/Um9GlrFHd63u1hqBGOJV1waDQ6yHaKthUHKjAS
lsMPiqhWBq+EVjhFfvI0gNLoVGi7F7UXNT9/Ur4zniTX6qrnwosP0ZGDBl9CRdsgMTJRFmCiL/Ut
PXbVy/VHJYZtO8s9kachBEyZEbve5Xprp3rh6l4v+4VTZNfxq87dPQRwbBRjBb7e6v5ZA8qWE+i+
Vv+WszFRxRBi8ejMy/omgGl+qzumDzdEaV9mXXva0KzaV4/os6gX3JRSCR2G7mgVGaFwZ/fkM8Yf
CKt+5UZkz8KPntHGqtNUpxqfqwtCoCq40CEUFVtSCsOqyLb7GIbUE3va4Ypmq8FMqISbqWEZi3m0
W720RkyVF2mQz7CS8vQnG0IIhvCAm+G/Q5HKofZAFK2JwRyNTsXIRqzwfSMQBj2vhKga20dmS6Sv
oQVYHQDe6FKzyx2vNtdHN2/kLyPomnN5Q2LM4FgNi7mD7eKW2A9ZPrq7QOOvbEJ2/koph++g7+OT
WUYE5560bXXfieUaiYRkBDTvkTrVUj776SXbxO1CJHOzsy+g7PJsGMY2vgtOKsv6F2ml1Bf4LUkW
Io2VTsRjGckZPOJfAAMXx1bj3m91vQj1HfltRGFMaCnLeQjxjiFMgY6l6q1R0kTDk/f11HJUamgE
gwRzRJF79hEmFpEokcMKh3gkIPfZsuglWbtevA+8W1dJ1dH2Vpv8NNzQ/CpCotw0KmuOV6S1TFZM
83wUE0FgQv24B7wQNE2SA25p4st05h1NLdadjJy1nhpd7pE6WkpHFyBAki/5NRFMNND5gET2/A7l
NuO8dGScTefzsIN5Gy6Z9iFBO8j0gHolKmVdZ8IXnxMyH69Gjp+BjLKLJtq1l5beLBSJ/nbL365O
R3jHn84zzqaAqoVd9XkoSTROSSs8uNYNBeh7r5AGmmY8kzZLmdnK0MZuyfpWNabKdAmJ7fQZuBPd
F7EJPftHBXipOu86A1Qzd/7pxxULSV0WdJin4GgBQyEc991qrhs/vd8OMADhXE6pCRZ9wi/ur9c1
xGq1EG+ritjQJLJFSNvkvLVbomF6YHwfcjFLYgkk63pS5sRBhvyJBkjjrWwdxFBhaOtrdV7gRi00
WP/K1N4g6AyaCPM9cQZkYkmAF62uAUlzFszlp+l9390wI1oNotSIdUN7HKStppiM5DrW31QowSMq
2dqsan3XtPBq57ZpLT2ADvXpnAJxKUdp5S4ynvFevYj2ce09/rky5hz8+g7f7pPFBzrZBsracCGR
RCJ+skGMbO+mTGx8N/a5OdJwXeTUS47P29pwbeertYw79B/V+30bPcR0vs8E9bkp8Ud5umNQ1V+B
162ebzS1ulz5v/4G0ZGliruiC4kmDDLzHlqUGdxAN14M4rRk0q7zTE3Mt7LyCjNJ2e0zZ5HlSW4m
SKo4FCaKt/+LF0LzWHzkrGzA5Y7fMzRNYeYzkOFJapmCy4qriXlnT16eG+r+h3q69bjWO9D/rcfK
eWRuaVe5a4LSK5NMNda0cfmThqpkWxUcyeFB9oBlhTSOpVadskHdUgQbtVU9kWtnVkvcrLtz/rVp
WG4E/OwHaWhclEbuag1CIQkDgS5/9+w65xyKL1UwsxiiHK6+Amnafx0mtm8+tjA8/SRoil63QXyo
2Y1xWYeo/5uG5xglRyd1O0n7M4JnF2/N8Y/ZF5wHd5x0MoH5QI6dQxA2A+tM1kPFni4HZxb33LGN
4XQ+Y6GsCdXMaenZNO53v7st6gnY+nsa1rzPbRbGVWfLPGkacRrO865aZ3I42ijeaPIBZAR7fmIQ
YqCHMJY3I5v3GW6e/Xg4O+ZyjglLHdKUVa0sxH0+I+bxBbPv42V1SWFtOfsADf2DoL6QfiIpFGx3
Gh6TEnxR5jGLTRZ1SzODLy2CzW6C1oxPqaC6/oeQM3JQlISvE7dC0uvIIIpEMbB9O5lUWmZTBxG/
CF3+ieDGRWs0bi4ZH+zqZHS36oRdznoqz+JyxmEIlAhm/NqVgiBB4YzAAGq+m83DuZYLuRTzVh61
YFI31T+jYuvfVu0AvOY5ZJBgR9tglVioeGY7Abt88L+6sb8iOZIvusQKDyqeASCyYYJYj7aB0BY5
l2ldEsX9OE2DkQBZJ/Hji0lQRotrKXNaXl+pF0MFPnLh/VyZb3iT+4Q4tGVaHn4bFMlvdpMOaHCD
GWumSQNR73GKR49gG1kyk5JUKD9fQeNK1CkPvtl5dBZHHdFRqP0Qf3Mgybv3xiBIrlvzQskTMG0h
7x4v8/wNKOLlMSsUi2ZUdmRtQ+ipgvmGKl1Gxp+MZWkc+HTNQSX8DLLkO/r+yaciuzR2XoaKVUM1
JqVVC0vV/BntbDxM4bp/5FVFbE8DtTKmznY244sq4GRr5dAgh1RIbImfCkkEjMI1I2dOzrhUQU3k
tIxnHI9shAuBbdR/KRRbd7BNiLlqvLzTYFfywASsvkAvdQ+ZGO3BiHQnpAifIaf0+7bE0fxbE6/1
TZYMBe1F6fOUql6nBbN2+KW0ZbZY2Ew9+fBm9tvUlSEajaRzbtpvAZ5y6XspOSh9U8ETimBs4Hcz
W0/XtWRwHW6rXwwOtfqfJpUWzg2SbWDcEc5qpvrCjqLquWQt5fnOXhCUSJ3RdPSI33ZqzXaCA4GQ
QecKP07adveTzJGAzj04fo1VCfJBEfxqxhidUdP2/aH9nrJfrFTRSJHiH0+B8bMHt40sjiPGY4ba
6P8AlpzVS906Nk6uOeTHMtLhPGOK6qFYp5aSjrTr0AXc8KTqfzkioS5Gg4DdTID0vnn8OFlYhwnh
n33413VK3AbgYiA99XA2wmYhKvC9iCqX+bijIXjFhQrbJMN4Kn/gjhgX3gcfnwlyNwrHVGwx0Au8
0ERxREXU+PVlPDmDT2dFFzM14DZDatpadT2fTfcAAh58PC82b6vP8syjgVG63t+4LoaWlChxx63x
GkD5SPwQac+i3wpcmCj9/ig2juONd2XgN5SkwQw0SohgOkm02KdcCAlZgA+Bi2aWXxfMaC/9+4qF
yQjT5WYrimTPVNSqGRI2Grgr5Ze+1idE+Q51i7Skaf5haKiccWhOhsmlZM3uf1FuXbMraI4xETr+
VBW8hl/sX6c6VP+CUE2LVN6g9J/FvqP+Qy+cwzWxUll2LKvkhb7e/yQM+fVgJR6XO7GLFxxsSMTp
i0v9MYNTAcmRaA8TEtMK285CzkHCgSQ0pivRq0bdmauYFJUz6bCymepV0L7iem3b2xpsyx985mhh
wX4tCc8+yCcNfC4AHmNY2BoBaz0l3B/Ixd6XLl5I2y44J5nDELHVRajXpvf1wspoiej+R+nGfdPC
2zMqr36eqPB3DDKcKmK05dyfsNRXB2yJpt15QK84iXAdH5YnaA6rjTm0H7pP2+l+4F8AtGjOc1q3
ouEg55ex2Bmap6mQr8zyqMu4Wr2Nz08JxZDJHkQmjDRu+VwVwIMFNdmpUZcsdR77m91UDblc4Kjr
b41gWJSAyVXjuiMn9kbJNd3NzJdOZJJm0TGNK5coGWCL6DPmDUBbuGTeGn0TXw4xjaO7DoVLYY37
sgStwMo2FrPUedqCh5lH3x1nsffw4PAYQILU4AjGz+cyCu+Z9snIYJxdygUEQwjYipRU/EMnKJVj
0c3IsI+bicT5SvpqPHnXcDeqYYCMMKNwlTjuziUIhtGXTt5rwWjhlrSeof6hJvXvR/5+EfW+6gXt
XH0EJXLCMSOfywqRrvJkzcYViXwn3H6JQk1QaTnO1SkYjI8fcI0OeDEmpGDeRxXGFCs39V0NzPG1
f3kG94rKg8bE6JbXDHa4B3Ev2zRNNBzwIoCK/Dhh83RLotn1cSIJvr9xWItHbVO50iayp/KsV4Al
MRHDslDGB2oPLN/IKvZv7GyUnUbZqqyHOg4604hvzQOE6zImyu00kl7qPlXlw1q6rviA0789fXAD
mQ1bkoPFhUSnySPy/CpfqyodDgMfZ112ZZ5PZWuublvQEXjidGPWHcdekO0nwjgXgzG+HCZPuRH4
I6PdJVQSpg+BDRw9rRoqwoEBCIWSdWL2vtS6Bjbnk/2Dw+DJsz4YdoSo4dcIg3oMckBT9/ag39pv
dDRtBIIPPIX0PUSZDV12F/U/CfkXN3rs/w6kZTJGxFAP+moF7KNVL+KkukW4VeHvymv2wl92fmA+
b6hP3OPt2B7wbHkBPYH7v8JhGXNIwKqrJn6neIi8N1mPPKX6WSZ2VXhcITeTM5aA8bYgCKbkyoul
s/dFpVUNJsyX/z44JtPMu0umofnGiUFiX2Nt5DwnDm6qcz9TGrQGPOUIudPmhmjoCX0f+cXEfBY1
KVcSy9+RQEFWtPKbfyMALzHC2on9bWkuaUpg9xZH0po8hGDSXuvaJZXY+OMUpP9gwmG1QY3Pxw3g
taMsUJNR9k/bJHRc3XWG0QYojadwdBIXPLpAhmtd8UU33fOcBu3J1+dMghBS2405YfDNn4V8TULs
4pAGnqFXBCMa4NqW/wcMEsiS/yRsIkQva9947Ijk1teMTN36K2Q8ePaes+RZSPWVDNz4b/lYdnjz
yqH6qIj8LKBa9foZ3zzSb3r1xSJOQqL6olRtTUqh8NfEEvSrmTXSTRB9KUrToGddxXPdTMBjYXif
hb2vzJ4q3yZl45KK6HSvycbJSYdh5xxwhjlMQ/CCtWWwaO30TJmTDoNxfykQmR8AeHujDzMVyrje
rJ2u96rb9Wc7KWAH7+Jc2njtc+MwJl0jVVzE9TIAraJx35rV+lorTIILW8F/kw7GcpDTVgsEekaM
0JGWh0TkjTcptDFb5037v607xgTykIqHLjf5ZOAB84Y4Vq1LWpmWq49GvpgW8rCVk6hdl9xyTpm3
HcBDh1evXsFXlAXF2MS0tMuRcAh1a97tEb+QGnayf8AnqeuVwdms6I+wfS+huCFq3TVQSWiTD9Rf
W98kimKm43wnVlxlLZWQRt8Mg6+sor0GtwakhXs2GVecMiLe4QHpiYmpd/jWDr+5RFYwYR2PjfzA
VBv4nOB8L+7k4RJGS8TzN5EjNgZ1eg7owasG8Yvh5OyfMMvrA5d/CKGNHqQDeudWX8yR7hgIv8c/
BdCDqtPlbVOdOLYsDHos4tQwfTNwdmLnneU7s33r6G+lNqxPkG9/whpEWsNhZyOCU8alFhdZNVoD
YXwji/InyxbTcA6QS8X1kz9EnFnWDwItSt+i4yyj0+vC4mXm+74fvW2YXiHEf72y0yoTvoJ3SobI
SNruyUwK/+yIi/5xrdlhI7BCnevIujTikk1cBALV1emwllHGTv91eCBEmWv4byd8IgdbJWdGTDOC
qb7dKOUQ6Tti4nR1XGBtrfyYeGUcBOBAAekE7ilmmyIl6rCw7fKTaCPxfxLQ/cVlKtnz8yYEzYlL
OkAx0afTTp1IiVTjTZ0a4nRyI6abq2VyDypty6tARPSmbkqsuaSXNLaj6WZnsYePtvU1WqvLf2iT
WhJwVTPXVqkJmXy3eBh+xcYM6WJB+iHyWTwcXEDCOOdjgWiK6y8eE4kUpKpxhuy4PKjjfFDHHpJR
iywdO/Mn05fx1Mf+fYWCTFZxHtHNWQaJG4p154E00hmkJi+yRS4LtJzZSei8VZ/+5wsthRASj/XG
MI7tHLw1UMJSUfBriBvea7StOSSprK0mABSavNhfgq7WRj6xyLpgN7NIVEyyrnFAuanyqGo+wBVe
1QvCDJR9FOXtwweL7IvQ7R6xa6K6DBvLQGrRm59pCAsCD5qFT/ReF2g/VEdlyTczMeMQpoeOsytF
KTfiwaDVa/AcivrzCwA+6le0HQRZkNvP0aNnhRNonJXlVYMSsJsC2EoHnkhCuiGSlq9a/Z2nbRQc
Bldn82Hm/iqc89zsCfjrGwA9BSN2Krfyhc+F58qRaUkTBZ9bJywpP33e1gPQ8gzNAdM/klQSBGRV
55P22P3mPx8L8/NcqHpifYGiWHfjvx5WQ59OHL3ok+tmeQMDzJb1cR8fjA3TA74fDim99q0tT3lf
3Ic1PVKsR8t8O7pL7D5cpWh6XAI8dAGVldeevxXhs1uOFl88cYGRiLE8zcsYwcmvHpKLmtIUsRi+
6UJgFsz8vZDXi+0fdu4mMTM/ehOAfqtyPgKvFPt98yVX+/0PO3C87rdskNsIwD0PW/bChQzIOZat
FkCEArva0bDjqGbNof0nkMIdlwwDsu577d1/lg8mLZ1LJIBgynrAMFSUXpHZDPDUmJV7+g3pLXuD
+Bhj7dodQuLMVdLOP070vdH8Rd4Std/caLNCW8AyRMmk8R5IcAKfQ4ww8JqchSZi8vvmcc9j6IXm
kEousD/WtfaTnjYVSIDfWWw+Muho7TdeIMPxdOFv+B7ppQX10Xxe9Bf1Ghf6TozKUYoN4OasB1yW
VFubTMc1qMsO+Pae+5CBIIc75HovrtJZJVtOrXC+uqi3C7CxWTKtHlnsMp/KrrLfEDmsYIviCXPn
ua9qgAGc4ICCpFFJ3IFk90Oi9Tn4u8GU7HpQXJ9X3H4RQfQLIrFLjFkUJxgTUopI03e4M6+XmYSf
WLxY5ZgradGSaOXP118PLADhjWdh+fZX5kbjaYXQyDXDG0pRnWfnR6jKY4XdlPmGT/bISKA6mEWh
BWphZ5HH/DNNJ5sH4r4tS1UnzXPvNJnpN0C6WHlqBIlh3dxox4/QDXW66xQXNMSQsjxEbCe78V3k
L9lOZFM5VkXsx9/0uYaigmThIO+P1ikBh16ZXHoirmAEyjH4col3TEDNrd5eUym/u1qaW+/fMB3H
udgordgstMjrmcr5D/0UiWMtMZq4vuZL/Om1hPDs66YcHkgrGEKYhAmQ6O/7LLW/PgAk213gMJjp
77uS2Z78RbtCJqCkx/t59mihknYmYrRaQhNK3IMJKUxnbr1w1YQ43yvCjQKMDQVVEkbqCbPmhBTM
nr3VSe3f5FIxnYDSFhFskFqXvG1Vmt8AOmr0tCy+ABxTMW7x04F/M/Jt+VkDRt853tO4mBxVRC9U
2M3r0l1LbYBC0l3UVPOaRmpZer7aHwkgNdUgk6k51AV/dV1PvYHDCzHXIG/VapliHJGPrfACwFKD
B0wbTxrJP3naq3HR3zdMnZBF+6hy5zymjZXdXSxzLjnZFWYUFPm53tO71r+jtbtM5S6Hm5efq5sj
sEvB6HbeYV3lvO9a+bzcKaVBxLj9azrcLn8TLq5M7e7ftTEluQt/TdLjByw/r5jIiuI7GxP1Z2Dw
hXQzATS61mG+wvQVGOKbtFXVWuyYUnW27tTEWfVnxRd1So6Ok1L/2C/tRNCyKzutmmwdzg3BoalH
WzjfnWdZ1fcaisrfwalRD9wqes4XBx3pMe9anoXHTfwYgIhd9sB88L6+zfOggDfsW1uoV6fu423P
ud55MJg3ozWIEg8wdmxNKQw5Ba9qYWtgDwX2XMTDNb9Q2oXIiwcWobYj50/5Olne9ZdzRH8svXvC
f/cxMeCbkv5gh3Gt6okfbdqQfkgvuyvxsNWBDgZI+rYfOZmTGyWmQpsog938snjH+kaIjr4oy7nw
y6ajakjNyM+HBHQdqh7mB73eypjdtTVUe9jb8jQ0WmJWlCSjD5Lqc2aRYonZkSDfrSVJpghxTe+e
UlDYqLQIiagB7zHoLa/WeH+8/r2reO0QijNJ4r/No7fivalOlgCwOwoQ6lOLVf9Q7r1kDDil92i7
usjNG+evbHgEv9d3Ge+D0Uwqca4z5RayrBkthAdyU2VlQ1+4BEWnmcpBCTPKltq0Mvz/SMATJdes
JkqoTkOYDIrpgZ8C7t/62s/LO+sF6fD+DyQ4j1Px4pGvxKrUh9y71IZ3SxN2XIW7GycfasnGz4/r
95xhExUUeRjAYf0Siq3zM3GzyB25EtDOJlosci7/32g+cJS46SzQELU2WUh5lX5haXCKUSF8Ekgh
ugHmaevEgUpWzE/EHkQRtKoma4IHk4hktE+VuNe0j5B4/+lqwx6gImOvkkabEEPW/T+Ue2gJNwCV
3DibAfCNvidy5pbzuShK8kSEmPi1ik7LXpZhIKLJkj3TNnAJU57Tr8zfZzS9ZTDhu5jYXPSQCuUq
O4jB/upPlLwmAMee5oWQT8YZy6jtUhsojFbAJN7Q7vT8pFttXrJSlq/6nNNSBsfjwAEYi94QlNQ5
j/YDW7bCmCRmXZ0UvBPE7sstvgBIoFs7r5vdgorbBUQEPIhHvlLubVFkyhBkDYIAWwHtxxhbl417
0a2Ud1zubtFDghc/sEghTQFgGsCHr+R2Bd9tmByTgQ9T8Mkepil+vzRCwUpQtPtal+Vg+mtwknhv
0u5kVYf3DhcEjZbioT4x0Jp4I2Xiq43SiHqij/Tvqjc1EaXH4n0zP1Fk/WfjR+BF3ORMsqFKWof1
OSj3jUsCWZCD2tiySahbQdcgvws2txzYe6g/2OvRs9gmZPBMjVuGQp2gx4LVXnJAPskX6o3Xpado
P2dfGicrN4kH93H+ydz5VMrdDDPtgs4erqeJCv9AsicX/9Yg9WkROvMLdiG2hYeAfTPn8z4qeyuY
Rp3ggo8SFV4TVO6JjI6WRbkUudXZuUiWsneSCFKUvGl+niCBHwV2mHnQms3z+6znrWigrNuLpnIl
sXMykdH74k6x52gzKnXFIkHRrv1nCSAiSPuARsRWGijOnR30D0IcLBmsqspM5yx+Zm9HHMsc3r0N
FlWg0cJMQLdLzafnZ5nlBzhUNYBnGZhBNlvfMNVSIUAv2h4CLzL49oqfX/XYHA4rbpDiKPccvEPG
2cOhUNnWE6p0nB4EOUzbOzSfkCLn7SjulFh7IhNlREQn/Gz73YqPioLDWQsOJ7+ApgRp9HohZtSY
8cZ0i3NYJRm8wuhANwh0gIb6+SgUkCoiGTYZr1RevRnVdQPj7cSLeiDCAqnjc6abLYAeUqGAcdpU
ksJquzPHX5eVFclpEV5jFT/NPIWOsTeQYAksfNGOc9qrDUkQY8HBpbmO/KpTlX6FQXb4nQjTgflz
0pPQuK2G1+74uUK+5qXmgWvn1EgALyp42fHK4OZ5rblE3lavf9AoNQMWxPo54d7tzZzwuc/uCW3z
mwH6pYDN97yd0Ae91N8UhKJHJnUE4Jk6pqjGyQpT1hMRYXTvTqZuTJCRJsbEf6udiJsAoVHJ0avz
7mpOx0bxoNV2Ah/erbCVKEmgyaiv6+WvuRKuoo53ajgjXNrII4rJgGlObGK5Q9c6cOFrI83hCjsu
dIk87taf8MpCp2N4f3I3ssVeYm/b/OM37MlszUkb7Yt6lM0M1Kwt6rQ7Pww9C8V7pAMgwcoQ1BAq
W59K/VopALtX+OZc6FIQ8wuH3LGo0iFx1XzVVYv7p9pTSwVqmtOHeUexOvbYahc+ZVvpt376sV6O
RkEK5eO4kkaehvjUZs8DAj08gApWCw4C2WR2tAnXOv4NbGJvj1MQ4NCZvxkPjrCYbR4Te8Ng9uPN
GInVxj6LQonr4cLyoYsGxE0YhvVrewiKmaHq97QV0zutCTpXD8qfDaP2l2dy1Ql/vU4fGqOqXKVm
Bg7n83NQWJMeOedn9mLb2XzNJeiie3E7jqnRnLAi+ieavo0tkZV5q6cwTHnF2d0eUn6+QJkP5gQL
cyyNY4w9hv8FVpvfwv4ATf2HK7fohqfn200UFuBi+IY4FHKSPiMCTekQ8n/ozvns9AlN3KuizDz9
dJ1HESYz/Cf4WdjzrO4M7H1cuCzj7ujc8XfPr13RXngbUhdSGHhvGy9VVgbp5aaUJq90jK04g02I
HOfPFs3s36HT2PGX41jzCafnuHWRLfOZgQSnUGxi/sglXXgrg3EKSSykqdrnZGRGIu2ayEaeJma9
9FUz2YDYmFUGx4ajx4io5sATcJqAPxOuMpf33bvcbqcveRqfkcQ5bQrxlT/c291xmJ0PekYtjg7t
sI3jFdtuMg5MrFtqrQd75TebAmKzVgaOEdfTghiatS7BxU5Kz6+XVVbCtsJVKqyZpkSy217WcEdo
g9lFCPQY/+q3Jl7nUp4mpZxruwRchBwEeSzfBw3booQ9s2QV+WfOf8yYsnSm2KyRyFsoH55NZvWs
OtePUEmad8AzhYK7xY170fpcJKz+1fU38Bh3TXb20/RAHvQ4xXOcoh4tAfM6XhDWrJ5hWI5yvKJA
kGTaOegqipqy3frvgokYqcg7foHr7SpfrZuAqYusYlR7MpP+/owlf98gYVb8AdegBHtJLKht/4o1
NkuH0N72ImZKSMP/5fARHswLtrZ0GAAv2eav7lJVKd/4u7axV1cWE7kGFlht2pxN3yM4QegUUrP7
y4Z0+ITmVLdbJ4bH9SEcBcE9SuQxn0C8sptAc51y2A5s4XT5NtUaJk3Pu7khEerzoUXj/5Y5b/pg
/oDvQnAAQgnhjGQ1DcOxbhDfWs5dtv8xY9svhy2t+NQ78qzJM66D1/LZEqGqYOt4WWKmPxh1FKh1
xLwuEa2qWTOXAVQCH4jMzVg3dKfX6QUALGMV1j7b3T5RZSjW0vWLryaw5ktiuAH0mbmFXvpC4beg
0Zymb33c54IJnpj3SdYSEPhv8rp6RKgkG5SIPnh041sooVrBSAhkO1O4AhIwXCikF082un2dLlOZ
K85VTbDK0Kxt6Z78KADphgzToB974NTkwh/LegtfiHFnhAvu6pQ2uHMAI9FZDjnTe1kWEpAHSUN6
KAPk1HcU1QLgFnYVCDIbSFoOSkb/NKw7UtLWzfVRvCjsAIS0XUqzhxKTeA5+1ZXyZt54W4Dkp/Cd
hqMdvEHXgyO/K7kqrhKqrbDNSlZm9XZT+EN6bob99nznRH+HPnkg7FLRgzZjGUzpSb28uEY0iPqJ
qGZSnSO2El9x0y988YnJGTTVCMsBIbe9gHAHG2kgVIE5YxtrwCADj5iyxg3HwZgNNv/Sxoprq/QE
mgk9XgcgSL2dy4CAj1kYQLQBIzljiGrLCPNr7IOsjqX8Jiut4g92HEAlJ1zQAzwSvQgdKiGx9kv7
HQCW6ECB5xaX1z1wfM1lStZvBq2wJcDCQ47P8FS2YkuCPwnPkoQY1yNd8JyeRWsdtZZN07hsbWO/
7Hhd4OehoAK21ABRCC/bpjZuxwbDQkvogR0B+Jhno0bpmoYNSbbiF721xAExtt3ck6KBDAGRzUhP
uS/JlB2D2bbo+RUgUjq7AkmCfIsdAWsYlZH3awsBBB1rxquNixs4kbzdD3NMK/CqlO2V4kLC2lY4
CLGx+VcgtwI48tSOM2jUr4pU1RWOyDAjwO2y2tWb4F1JO8H8lD/kQBI1et1tEIzTfEepLyXx7rKZ
NjqPRMf6L8E/6la5xgEq3xwCj24q812SNWSD67XTQC4wcUvQiF/vgRZor7Mfxxzpzvo3zj5msyjp
L2Tv7RZQtUmEJI9EadeShnPEetuDZn15zuknED2Fj93Y8fuGm/kerFB0fPZQrNUWPvDYHdCVi8mm
9o58XmUvpMlUT8bJCUscYkDjxYUZ4JCGM9NLpeBHZeHvXIWt39LNIxzlv0/Sem9IaH7kY5L+OyPm
lNQGPiuHeMJ2G3G+frIjOC2A0Vzat6Lxks1yAila1pAGw/PAT3gmhRA0Smpet6zz6soMTqa5XHJG
EBLxCdYpkqpdKPOwP0OuHDmqtl3bb6Hx+MEd8NO/Pfnqqj+9upRdWyi/jaJLJKEv+FqC1OL5JuTS
xrbNR1A7Mh0eDLWRfAVGBHEIB/WkVnZ+mF/XLfMwodSes7huX488xUweTNWh9OhqncPjL3mi80eE
VeAf86O6cvkB0/lJDQWzOPRyNfGBunNaicfhjMqLWWbr6UQTCBBCh9LmKITkKHDdFyyfpMfKF7CJ
qdzTulz+haTWfHFcADPvpCsuOHFnfcqRl0G8nTYgKME4vYioYkIbXuY8HBlccnfPTQ8oT2MtfFGP
7RGb/DTT9w/g7OC6S5WaVocLy6enEJDsEoMosm9kPy7dkJy8zsViUD0UI0cYl2jmzVhNCDzWcApN
gtJgF8ATRIVO6fzQCiSbLb7ubOgZ8comDXnCCpBBS0glvMJvEfbu9/MdbJOkdsrDEsyP4qr5G8DR
wIPNLpx01gniYDBHsQRr27Z0d4XjfRhljnRpGGtDoiSZPGcJd6+RvHzN6Dkmpa94pi63idqcLzbb
CIxpTgoYwp1T9vJzw0xFog/l3tmWCIk4/obPgNcPHfXtXjTpOMwR8kb9nPoHKmK4/tgw+u2aFTVo
JyH6jHJ4w+UJcHJD+dp3h/Jv5YIQ/RwhQNs87+Vhah56lb6zp7yFaVzrnw7Nu8KNScEQmK55o056
TTFKEIu48xKHxpa8OfRvrKno90ZvcoCYZcydU3bSVuMV9JCH1fYS7uLhjh3h+MZ9EpyKEyr4+ltO
2nzChRLiClmHndg8RK7KHVKYJ2IfUEUrMojFd/M8PSZQOfGZAX0N2VA6RH0+hapV64JMK+S7uebS
Tegr5Tn142Hrhl5j2UIozAsOoPh+mS53flXHQ0TiTmZ5Sm1HflH610gnl/kUIqv/5IwXmB8wpedx
s8Ia6YStlgZOKZio3+AN/Vuoruk8anpHo5ECKrmAyDi10vJ6FISHckmJu5qcrTMn6tgkq9IZd7RZ
hSL4d0KpEH2b0I/kupfE8eWsQT6BAwLewLXsmrqxNWK8gO3hLE7Rn0J6L9I3RuBndJNt8Z/S+jei
dTASAsDN/qAGws6J6g1AhTDfIQx1e7jSKswb9NuHLTdgE8Wx0ml2TJrX4zXO+fJY2+Unv7PpgSU9
j0aYzdvydm38B7bo4FwhvUiDG3dt+6t14gwh/Ooa3oTUSKnJT21lLS1nzNassdsvihdNbENKdohB
xXU6Q7wwWBchF5vpE/aj6kdNbFLgJc3DO5hK8oK4/CBXAXDTKEDb2ytfUPw4EUNNcbUYUHibKnB4
m/Xv1mEFt+LDlpmdgmuiMPc8c6FtU0mIEnG72javFmZ+zATVUaMGKTTtjBXBzZmCU6gADMWA3nSj
4VMmN7dsQ0Q5bVi9hvQdq90Os3qmPj0FLlLadbLoiXqIAMeuQA9079ckmhIZIEe39ZbEPSEGrnzC
Khvj5ErDnOS5Q/Lex0Zecm3+u0eCGSYqnkeBARF1nprbMdMozmmyJjveE1O+Bvs3JvIzD0mX+HPq
EM+bLKeVEx+b7cy4heeGpSmYVDmBYdIZ0VuqKFkHtnQEvcmbWssNafylXwMkggifIXlc1COwCAYe
+omMHiX0SGhrW1+mw0WYOdtOaiXgYE5P/15q8gd+VLVe+bFPLmaMksSdTQ0jRL91JERsMIZcQUOf
aEhW/GgOsL2cN9gRUOg/cjTENeZ5xSlFrO8JBuVhiqUkedOSYySKkRlKZJq31YMakfBSi9v1B4H+
hHhrxJ8tgszba+RENxNPLy7qOwsz0bxD0Wc9T8wFbOlRSUdPUfvroZtgFOt7PODfdi7wKJT5ROxy
+5N4y5he7umppSqIrpeXcxcI04dnC7PyjK21xnF0IRDBvlRwtyGPk3HiKCUQNXsCcM70RbgPhvT8
8IPeddCDh7BF+YkpPTat4RFpVwDojnYtUr2Hs0QIcRpOvLdplZEO1e2BgMe2Gw8UmA/VfR4FQ+5R
DPXDb+mDZWxT3XcLGXouGnUbaCurzL8Sq9cG3UgDxPgKqNDbu9zNTIBCk5BwsenpLLjQ5tJL01bX
0Rp95fWno6hV23U2SNM2Zya8MnzB/5wNTBtLvAuq4mg+4drNaKdyUjIljYG5lyCUpjbwF4+agh8S
9Ohx8lVBf3hWeynktAh1HXI15vs0fQUc4yq9IXMGrn3O0/HLM7WPaidzgqKWmtH6jwVM9o+F4WsP
+jtGn9sRqaKI2Q9Ze9BJ3O0lvZeqsxeyhgrIMZBsV6U3rV+dEuSr1g8TkztbVj7NKQwgh4UWw/e6
UTWTdApyPMJ7qgqloARV33CYxIcd9j4X2jqL6wnbwCDSjv1DZNS0tMv1yCMQMCzaHse7gDEu7x3J
UyXoJkCGlB4ElVt+qiLZbx3mGM8IGTY3QM9QRwy9vuGLTSzh9vrCCOP+nqWTkmSmkJ6lF3RJ1T28
K4VHkLrKI0bOTRze2OBuRJMBko0j2nsVtAEVV286CUSDRoY/xJ7vu5bIKE4YeXE4qXbkr6Pb0mHW
oNQ4OTbO2Y8/EUYWq9AJzH9ar88KjLHM0//KfIFWOcyVff0h15s8iDmNr7qkU0/kKlRUjaT4OEjJ
IVAyxIGdNPcNODkR+NK5xpURhJ5EUx5e9PXuBISpb2twJyiNCglCBgFONl6EvU6xM7oyG3G9V8vz
HPrvEgVt2mxQSWrew+02zOHzo7QokXlXRLS2rlLCoFEi0+EODtBhbsEorF9FW7jKS78rZJrsAvLK
CI1UbHzC7iLu2Tqf8tIpLyl3hskwgkFUhzV9NvpI5HH5FW/e93xJa5DyxgJZXMaeOA8bWXIBrEAS
jpEBQ+qEbOwabIGKz11SO86IAwhA9S6CRPYrcV8VWnZ/C2MlceH/uRqhKZXPTDRWoOunn2DEWRDa
cpJpM4uj0UDTy+JnPeDniQUGn+l/KDRyXxYURFlh3SU4s3lkTG5ZU+1mP2wsZJXhYTWgCsFTa6za
ltbvpgPAzONgfyN6DGWerSLcrpcNaWP0ZhsnTcAv8oOkipDJW3H0lcqmngxt0la3qtY4m1JcPnIS
g8OXK4bHwWdXw6r3svZlNxBaTWAiJYiEbszoAcMyrQ6tfb9gZCM+xf4ThrxfobM7KI4v0H6nxRmB
AIpMDTr5id8eE+BPxu76ywrqiZSgPt3NMgRN4NuVREOB0Plm7clnc7UHs8kxj+BRB/SffTpM3xGl
A9hcXj5iZbf2lJHY+KQqDe+z/2QDfmVkTsIpHgry0vb4ltty37o4XNwXTILUt0lVC3XboqE+tQj+
phB/Oeuakjtl1kArPygXhrDLxJot2dyTU1yetvESIC4WoEbsAQGVxzog9FF0FneSlz03d/qnnIIb
J3IYGUyc1FuiiWFSHkLZj3VNhN8x9SDXbJdX9/OSp9Sqs0YlQvzoewA/EPBEHvkaXPZMgWyv5Zgr
i/xYgNybobdBUe3e5TVPY/MsQSdxWG4OzObHdUnc0XA5lPvBXSBPTJymNZrdaVN9ZVZGAtcsFEnF
PVzKVsVMpHlXaIE7qUVfQ8NBWnFooD7lu5ejoqMOM+P1/vu8ZBOg7uCm8+BOYwVU03VF8GmzXmv2
iS6qzQ+3ug0F1CTQrShCKD5+PpJ1D4z5fPdEUGxDqMEnpvCZtftTP28aqdKYKJNnS2QH8IHyLROw
tYyWL0BS1mQM0jfSuo9cyRCl9zLuUGE567GzChOyGCCLyERP6iFt71CZ1HH2Nh3RFN1cv/zNEs1o
kDMPLK1T5X/ArsHyk+Oxh0FWBeGLxjvYQH1G9iySUJE0gG5Ddx8gZlIJjv00Q0MkwNUoX/F2i7hz
ifMUnYNbFqRnOxh3wizXvVV3jS+LpoPZAkdaTp3pj7EICPbpXBp32B8VtSaVCrSkN6KJC+y4g8/2
ExBWRuUTpwhpp9bsVWMVYqslvwtqsivbyXwhxFpttVNuCVZ82Wc4nu9nHveVoCwmVzh0Qae4Z01W
X+xobC10bfPsdOGktMdZU1uho3drRKgFA1lglPHRmABM/ej3ssdzwJL7oBLJ8VTxBtME96SLkn8k
3BJ4xm/jxfbuqrm7+SzfWqgeymgG4AmzUVXYy8kIzuRXk5IThu/XQTYh65j2UpKfMQzl+0ogm4ZE
+Y6zOsRrOCtipAEfgbOhff3rEYVuiFju6vDkJktZESwqmedxfMnf21R6UCO7LVxfUQGF+RHag8G+
jgxqWVRZhVAq4aM7zQfLq8p959I3dLyh29zIj4xQRu3C/fE1dWaqwhxICRTNBz1J/ja8TxALaB/M
WE5tDKKV2Ao0TJmmJO1J+2+Rj5VJnsSFdPxreQVMvVJHC+fWg7T/fJGGsr9116jrnjGlUAmP/S0B
xlzNk4Ju6rdKaNN0kVPlpg+Ov6uU344RBo9kxTZ19iOHqdlI8boz84I3rGo850xIcOA0UNREoO92
6fOTMR3f/kQ4DbTf6DfxTWud66L9gi9v5srQZdhNAHo9v4vEexnC7HowzUqwvK2fdeldscPAUuFu
0X3wfHhwJb9CIxxKhcyRVJOyxS8CuMT1T5A/dpmpqDHgo95TDH8amECWSossA6LsJHiWXbzMzdnt
8TaTJKf8gBcl2NdDF3dZP/0CjrqhVAzosQOj4lMEiIsS2UV+obCpltLfF84C02mbH03Bdg+ohJzt
Qirz52X8OGu3vZ57of++9Quj++x0GUY1fh+tvg9EhoHthTcJ90vxI2Pt6pa7eoMtUHBYL+XJWtJx
rsQxb7wAkZb1BZNy/V5aZ0h1IjNbnKzxsB0PM4NDDa1wJga5kvgxdRQajFPi+oA41zk1xjIBVuBs
vu3rBHy+N2P9QkQwcZ5qPFHZIn/okCasjZlTCepSxvG0/umTd0KgFVLps8QJpjEgKSIGkuYNVFu4
8EqXDDnV2R3xaHUVUTUPx+ujVSWW3WLBNttotUxUJMKayNoRk1RucrohqAgXf8FcJQJ33fbe+bBG
FE4d2r5LmOEX4nj7ReOntK4nQm0odz1zRNPuZg7DggRFjijvvvw+yga204UtEWQT5bn4BPob5I5n
dCK8L6f5J64fGDljtnq6QpV+6sOTVwCM2q2CttZdvOelwnegfM0gSe4RcxhlvcD9hzpQiQfAfKXZ
mts+FL//vs+sR8LI7n/VGqwu7Kf8xbk9DsKIn2pN7xYwlsFqnYUlIWooRTbMnuG5mr2qPqt4hDmr
2qq9ijA7HZqYCwoqBxTcYdM1kGJHvTMPnOcHXbmDRTiCVrJF0QdsVSoR0ZasiQMozUA7qf8ZMp++
yqf4zwkRJqlh9wWjNBHr14Cjvw2YjALs5T/vEXaWhSS5D1q/x9vpG57gz7/sVIXkMBk+BhMgDg9x
TS/nGr/gnXXMCrnd0MfvjnQipaONEh8vNpWotNIgDfQn8SBbPj3qNivN6Rjm3BxgRiYHue6kBjyr
MwaY3nxWRvMUyry2XvnYgAT2R2zWG/Ew8P0PJHAXyjMAnJuE1jynDZrMrV0K4re8C2Mmsrd/mElA
Nv2XbXtKY88r5qgMUjgQ2d3FLGHLYUnIt2/aMeIi27h/YAgKrqgn+NM/H/PY2fiuetLPhUpz3Qaq
WAP6fHK3O//uEH0RQRpPBPVZOU4aCVBSYG46/Qm4wrYLKGDECSbmw7GPXT7tvtE8yTWajWZXQn0p
4lY0UVE+SvMc6qThmx1Xr5odUKEVqlVBNYzI++hNNFO8JRd4yQzoyNv4UcHTd0KaI/5hWCY9Akwz
H6cMtRdoufnALTo1J8PDtaeJBofElloCT7y27yFQ7jQABZe3KH0wSKRz9I7wx5Ojz2nnns8kPxAX
ByBvvdG2VpbLh0IRnhbWrIEoHXBSeOs8IK/nBEQwU7YAQmrVJOQU5ocxVP4KnpZzYXkLuvtIxiFZ
wVOHbIrFkv+Q1ODYgFMU+MGe3sodlL3axvIqGvRkHbKndgfjGemGa2y4B1x1McDO+aBip0fe7/sK
moW88QyVvGQW8BfKhKJyY5frIPgUxJg1WRYvIu1Rrozu8ikFFOzUITpv24Y3yi8yvhN/KKBQQPpY
HVKbFq+va+qOBFMCsC6ykg9yGdKDEBRnRoa0funws3EVo6EdFNup48/GjsThV1GyFG8XAl5xrnh8
ev/h+QAex5c5ZQe/cZ2LTY/9LscgMixP/ZQQUOC4yzdmrXEjnu0dfshTEalQUv0CzsLBfHQS31ol
X6KxGwCx212hvjZzwHILcWAaHfBZ/8CGlZd5ADLSChyw7xY9thVP0SMrSeHrn8YvsxT1vJ76pBW2
UkZjusn0bKtgUb6tRMCf6dYx7yOs+cbaHF0/FFK7u4vulvF0WqQneBgZWYhECt4Z1PQ14+TptB/E
cFa0ye4xgAI1uhc+QfuM3VBcPWjj2gpmlNX6T5VOSSB0NkJGru/BCGdlx8HxEDJ8pzad5/WKuAi8
BmswfeIR+BK9BScq4CaRk+2gULOzkHgFFdgnhdyJtasfHUR1uEd+wcwDIB6Xypsm7Tpuye9igUjU
8oRc9XcnqfhxEX/Zvq1K3ssU8h+C3TW8DNfQ+2G1+g4sdeoGKt/RWNFhdXvs6L5GsE8qfkQ19+rv
HMUgdfcD+s28VrzNJcrvacyXoT8cwsfWQuzOPkpoeYSv/l2YzpR/SzMItvWEjQrz/U/HtRFJP2zT
xAAa7Le7rn7fZKjjsZk4Zj+3a2RwFZtUUQRjSOZGaX3nHvKTch1rEaEL1jfogEzi7S98CwbRuru4
kGutbG29Kpl63ueYlO70LNpxHKVt4GkGyXWtrK6jpHzr4j4iTbqsG32xo9Wb1tCGymlzWFrdzD9x
oYvnv1K/VfGuDJD+DktLuVlDIJICOUkleJn+kCPu57noiVHKVrzLNcUo/lQ3CCy5IsWrUnebaYs2
OwYbpTw6kCkcb9bLqMXapfz1cJoyPc82IpZ3ZLFVGGQNyNaZOiCfbAi228B2FgEPVbgtl6ncwwFm
qAEnuNKdcKZmoPJ6mKiEh5aAB30Cy8BF19qTKFTvEP8fsFahnPOoBArXzFVX4E5wayeVNs07myLH
A2TPxD83fT9L6+hBUSNX/YqRmChgl0Nh+2n4oZHjFlMFpOFBs/tDuesuKwbkGfL3EhJDtaWUhCvr
u5wfbuPQ0voyAWhstioxak0bb2lF43Ugj7SK8uW0S0HadZGgnN5OwJ+kQ92T9Ftga/h/y5wq5Eml
GGpSdiNQDHPY0KWAC66E3jUmAFYK296f5MnrwiMxKCnmqA9i9ugXJioi7hrCht8gtzNsWzJDKmFa
hGdPMK5+q4e47gHsQ+slgZywfpFHkyy+DmO/orS2qD+TSUf+ljuLOt5hggs+tJM4BFOSeInkZ13M
mxH7BjZ3UnPczL9V3G9PjGMUPSPIuN0VwI7CgajNEq6evEAXYUurq+2SKFKE2t0Z/J8cUqNqHFDP
JRMaWQcxuQN403zLqO9H6NircbxNcy/deKwKKqR/FI11WzbjFHHjg77r7v+JMS00dpXQypacHnP5
k13GL27UejIyYpXDsHVn/Pv98JkSBOLTHfhsJwbpWMDrNxgyGpVnu7ZgLhqlnP03hLyQI3DnDRzk
l6M1Iq+QGSutb+YTMHmhmqfOK9g7YQiSBXftEjwIoWE3YZIA2dWPPWgMHkTrK8abnxL88Ern4XHV
KoSG29TWPJYI9rSujXmoH+nlbmJ5MnwRO+GhwnHJJPmOQDOB0q/+nlHESs/EYaRknLkI3a/QIIJp
1lPP46vZn8FLG/yzepTlx4FzuwGtQPiHTwkZjmTq1Fc31JKPo2v6tmv/Ha/n9CPIolL5AvgRTISM
eSxXH8oXfhmncDtHk2MMkgJGmdU2T/BofChhAuKyvZoXK/hIdxmMtwPuZ9yNBwQtevTIEtVRaGMj
FoM5IsTGgZ6flldPHTsK8mipUo/vq6SvLzYMOqvEy3m0M9OpIcOvJYO6vSXO8E9Ma4EbkA3bDZ1a
7gByg/viNfynBkrk9JKuZG2/0WywaqfuFxMbSHVSU+PnbCai7DjlpIbNkFvt9oQzNvK/cRWahWd5
eOLg18LsoMD5/Y470ndrYUfD1EOsZZ+qD7QpcnTl1+CoN4ivRQ5hDJgF1/N6/JUep0s8Pks1+0hB
t6prPhqXMydmMR8k9SgesgY+Q5FBQmCXlGnxM0LV0I0MVIp49hvT/7LXJLhXy+IOvd3WUC0RoL+i
D+ZKHrjDc9q96IIfHO8eA8BGhVGoBNTpUZaoE2zGGrZPzlC2nvDqrYOQixm+h0cJtOFLr+MiXZJC
gukSQmHV6AZ0AOko05g/ijnC3/4u419+gqMmhJ4lXD8Bw426C2I9qlaE5Ld0qQ6oHQwRVjZ/fcIE
dHZGMKBriNIuOmZcc/j3cPH7b/+xaOHyE7SPXekmi37z+4tZwi04eHEC5iL15DKq4PeUbg7U2koy
HNxqN+mm685kGPIQSLISPlJU28RlCTlL+eAAbKNZZVtxZygvgMRV0M3renSDOZmbj1YnDX1tYGpi
5hl4NzfnNEo+AK6J1aXZ6pUjHqEVjihsEorHwxuQssC8BL0fCDW2knoQ2CAu0oGbfwxiNFYjqsTp
1X5kV7uJuCy2Xat8eWwmTOWD3cDpQ3hWAr9e8CmBqPwjkiOX38ePcgMA/3BaCVTXFApmTPC8OJR1
N8eMV+flmHdBVMEz6nX/tHhI5IuoKjtk1h/6wQnddNrpMx9fAMEMQV4jKHEpm4GbG7hSKZgEUK28
0opt/c4jyqkMGMv4OTfYKKlEjb2ceqqkSg9SpfJMVCOuGr53JmVgquGxEaMFcuqw0VUATf4nQoPp
aEomDoSFzGmP42SO5SmJha+oi8o1D/57kwOZCQwPvUVUqishK19aOp/gGy0oydKS6Lb9cYzHP23D
2wAGTmK2/pZg/OXIlayXByindF3yJRaeLVZE/IuaJrN1XD0tsqHyfI7AWINw/QatTVIsT/KXMhlK
LR5ZN5aq9KipJbbCxng4tiZ9fXwpiCfsUHL5o1W2SQCz0MZ5Ux7+Rq9BEukMtCfW1Fp3kcwhmjGb
iloFk/lYNQXzMVeF7WRal3aHq98DgJkQRgohZT42GcglLK1YmN9Nh1AJ+nHFkvgNV5UB70jIOB0X
OvzknIldUa9xNezyVftGXINLo9gE4QqZCjQQHZU7ed7tToCEsFRzMJ0k0PdFVHfuAREkKExFZs19
VUc1b1YeGZAajaADz/7wc2GD9q8A4N0Fwtz0YAyG/yMp0RdA8fuAnR9S8dSr9o/gNu5ZPGAuGrzO
ViBIWqugsGBTGEqeepRjBo0F9bw9zK3Rxr1/IqD6IkuAW4hJFYBygJ+aswa/Oa94/SsIVikrUQrQ
Y4+boeO7g20uNVGqRmoQSIgL08vayhBH8wX1clg7IaqOsnZqB5IYNu/rR4iRFGf4ewFoDp1rBdO2
XCnovr5PmZBlamQ8kY7+ncC0JwT3zHsTU9Va7+0tEJPVYw0CdasxH67iHLZwPqi48QnkUg6IoYp3
RssGVlQ3zCrohGe+QdrAPcl+e/NGpAamY1fYXXE9y8G6thnresY01S9uuN1pP2i7EmuKLuoVRZvS
X399Ws54XL2IWJQSLIOX6DXBOqxnzwK7WVMMiYTEboqrbhFoP6V3Mks/m7aFQH11l/byvyR3B18L
j6zoKbD8SrpWYXqngtXFn2PP1QGgAvf7y+gyyQtEAHwD5UHIpKf5HV78mpuj+ZvFTtPv43Pov5XY
VmCID0psNCc9Kuz1BxAr9PuDSUmYDFSgw1guXzlgFSR1rY4rIqArS3hWdvjNoZuw6BrAa8D9Ucba
CA+4KkSYaCS53CXH5PO8a3dFoFnrgJAvuxJxiF5WOvSIpacm3JF59ZQOzHzoP7IiR8E/8MVBQ/1C
H9/TLRddSiiKhd7/3wJzkQuSM/fqzeod4O//4cjNSHBhXUumCsZAUdEpbSc11teK4yBihy1cWJIf
AI7g9ChQBXr5vNFXvUjyhVBEoe4ByPnu+P4MYpvnIEkWNFx0DWcUuIHm1eaLJJD5xFionlAnYREm
rSVRRGlugfWdyVQSdAyd+bbfIkyWQ4ipLNGaYUuC9yHGiYUKRbd5mw6MtAL+pmP7JchSwe9/uuwB
/5y4ZXYlYgQqQSy0LCljwdey94S+uUdEBz0G2blLSHt+MNcIB7lZX/utm8P0n/LT5auUYkHrpC3n
TlANrVVlRJvGiWTXeZcaeazGH4ALOkAyw+gLsvUgmiKo5zu2Gt1u3E3+xc7C9xs4AcYseXu7cTVW
zLu7NEzZjgwnzoWLqXoFAi5QLY3XZPAF6N6S/abtotPWibZDIARcxtR02KKeQYmBaw93U4kyfyKI
81E2i2TFokXCaCpuxdCCZvHrmyhRispsQQW+6Vt/KpeL/wNFYegsB70RrEQBapURj6ynIHWbjgEc
54zF2WpHq3cyLzMmKlcapKhmPUhLA+/BkBGRM2jTdTBiKpFSszVJ53cJUrKcRmxkdQvUwZAb31hd
wLQZ4bhpQZE0vdvke2Ga9kewBtLm//8+77qzFOJpiR2W45vRYewxZxonnElqusdIBKbtegwQAHIY
35VvvNyYh2nLLY2AoEasb3Hi2R9aOR+WxSE9w8t4xCD+12FanuaOkKLk0z/GuvkIr3PZSrged7rN
xJ/b/x7wX/vrmEOUNmayFzbQxyILY4Nk6L5MK0FCFNtzjWY7g8SjJfxh/+U5CegA4FzP72OEiF8O
cg6ze8NSs1unIUhY5V14Qur4sjNSQQtj9QKRsgwY7EYVR7bd/0iuSb3zfiTMgga+rhYIdjwiikdG
5ey7smxO7AFcAZrDfYoJIrtsxix77cPE8/oy22/EGPJPHjq6s8j9txJUY4HAzmhpkes7uvJjCc1e
eadbkIrmNqIr0TL3VOxMRzXZkarkFToy6ILnHChkHz9M97RWEYxSMhFFbs4ldaBJ0z1NqfmrWOPG
/RqPU15HYZkL9gzfElZbu/qw3sCWkPmlXK22qC8BJxMILq7/3bdq5j99p7WqIjtPQYE1uJdvgcWV
2Lw3wd6hBZSXUk0LiWy3HfeBw+/OcCErgYIBJUcu1yQUVY/hlF9AO29AoEPD7K26h+MxcDRFF6Kt
t4EMHTG8kL57+31KJ2qQo14S8ufEuMix8aHIuAOBRzPLqVe3PdGzgRpBDnxhj9F3WuiImIxnOMFv
LL6Lb1922onpZHFvN9OT7r/Yt+v33OZsm8KHqvDI2ISjZFLeZ+TokOoxVC9qGOjS8ytP9nOHedGs
VmpYehLaIszCDGfxx1o2xa0jUh4JLbNB7Hj1QYqlHTJ66OrcsPNtJasXAbZYHctdWMWVfZRhvQn0
UypoAYF5ZIqxBKQGmSDrlbeI8/tEIFMLFKMTd+T6PS8aW8uVoafgi9AZBThHPqRlVfU101I31C/l
dnMlnmoGCmrahvXJfYDrnDb9siCBr0F/ovgDGEOFNqBba+faXAf8u+MA1Zw/l5UDooJ6SSLBO0lF
96+5M8OBslE723u/pPZD34WL+yiifITXBjhomw1MWE8839b8EJCnOqT0a3mEIlYttT/tOb7Tnmsw
Nvdko72eOxzjWUhmMXe95RYVZ8pnulfyykCVxnMfxM5im+M7nNBU4VZg4tyjLewu5Qp7W+Gs+Go3
c+eIgDFtx5qbIVguTKPyOMerFGYw4gVO33N84vVFwHNsF3ezgSb7AcwkHUIenfJSyK/jGCQCJf8D
rljUmtl/HuM01SUBO7QsdatQHE8ybnCLo1MAvBY7QFbXYxRaOXI1I8gIgf4Reu1uTYuq8iFmApEW
/XU3tnhqH7TS9EE06mo99hOQr9iDAUVHlH+MnD1c+gjgtcGDosNprTBm5LlpSjIXKYKhAFYKFdEa
iDZakosQ6oNffnFWePCVd+Rmh9TgFFaiTR7DjsofGsky92MiRxW0qfIfR4I6I9IBcIVxjT1V7A1J
pive+wZF9QCVVxw8lnd/6DeQtSXHhNNB8Af2jasLsWGIuHMR+MkrhjIUJOkQA6bGUx5zFaT/IOC1
Qd0oQVZGwCZCtg3avMZxzCFXTN/RgRh8q2JE8BkEtFJ4WPsWFm37dnxYUetmuGnhV9YRK8ceIky4
4nxiWkeqkrgMNmtzfDwo9bpDXtZDzSZJWpvB3J1bZBfx0ft9DXNqOXwSUf1Ajl8RtHIKBUi82yDI
BkVvLsgkeHDFU9S2UReZGPvX5kD1daDENquCHsNirO0HESEUZQLgw/cmsUBTiKbwBA/VuQq/Eu+h
yunQuEi0pctdvYmJjrhfNWhZjE95xQI0uQYN9LOJoLL93cGJVOlBmN7gXucFHV+vQH2xH/9NoWD4
CExg3QMugirJA3dNYS1xTY3eE6lj3ae2peJbbJFWALmNcoUpE3ZWO35hsBDAKg9rv7NQwKJ8mBNq
CqNRZ6hVmAzPt1iBZsvwDLsideYulJ3uLlXam8bXby7yQwC4uSpig2OHYGEb9M+2DrIM2ccwzn+b
ZkvNUPYzOGbR16FujFzdG72zDwEer29PDHOTpi3tZQAiTQNQaeF7K3VVXJE3vaFgroGMfTnNu59+
RZJsBYCk57CZ/3qYzB6g7Umyy1IURYHTgV/aJgqgO93JULiyGzfH02cj/xmg2gSihoVEYJBEBTOp
/WJlx7A2ryhE3htyeNc0aFyH147DjZ1SjHKaLBJzYcYcDpMLbnF5gPdh6/SB0TnhEXDAN/hl3xZS
VsB1CwonToNY1XJkXQaUE71ndC1GBEel84+rR91GwJMlagf0gUc1JO/+odpmWYCHUPlz9HJtHj51
3gSl8yOqfOeKvK54PyhdLtxJlkRGml5Xj1ISwf2UEs2Fm259vsnZp3AoIHDujictq2bLXiX+F1db
V+wnFSq+lC3UaRmzdd2/RUmQbbiFpHr7IWfgL4xHDfqSmbhLejm12zQxCLT1pMIqbavB0trjlelO
o3H88LHT42U9ZXGV2ct2IGFIqTYIU8hU30nxadDPfAKu+HulG9QlrA/qiUseWv4NvDXurnXoQPVM
zFYyDO6yq9bIf66s2KXTJjk/zvPhJlJ9PDpe2nA2tXngJaa3Mjj7o9kqzCEMWz3DalZKgGNPRjoV
xvr+XF0ZD+GahunJ09IYxeHhHgDrG291Cl2j8qMQDAFnKcHfsbp/gPvNgtLfPBNXNJpDyDacigG1
S+evgTP0mDHgyCrM+/HjsSBkV3WrOV7dEAtHfUmjVw1Y56x6r4gK1Hsd4qCuPCPiy+U9axBJY2wU
rQ7uvSBj4Mcyz16llIOBuRVuGEAE0EW8uDj/DM1y2WgaV6LOny5M1bJxSGXThnxr7kIChLXTxpNR
z/o7WN0eCnOm54m9JpqL1W6OVM+uFJw2Dvlt+n70tSXyD7pGaOVN9XNrBOk8FEoVL5juf9LIeKuz
V8EY7u3XThd8Q++VQG9vqHDiVALxZHpypmFj+vuD9rMnPHbvzU8UVNpBtteykKcdi523Dv3tS9QX
wF++/+pyf1LOGtr6BNjitd/aqpI97uXX9CaulpvMAkFSDMtElMYRtxSFLeOpJuL8Q+rsMP0kXHlX
u9lMz9NuEzYBreOvd7UuIcX/S/F0l7RnwcZBB32HrIF8aQF0l/qJju8s3BHxeVkrz7R/B3cyrPYH
iyZlExPzKimcvfABrewpqWg7zk1dsX4v/0nB7zeD1vH3co8BK2tgAPtCjzy0mHRsWWMl1EQa0bDy
jT2TqX1JZQSPGAV0fMfnMlgeGlnVQLThN575oBm9L+kC+PHz4LA2FtHLjnnbcYyA/tIKDGsXGG5s
EgzjdHPStTkoyA2b7dQxm14e+hIm1kFKQMsDcDD6FqomqLkvNMnYHn+4S7a+Ya0erzaFlGVRmw6u
AW+4VfES+w0jP499tWqfuM7bfCY1SEUZtUA7BwaV3HRIeNu/kOu7Lw7+5z1fqXx0f9aAEuaxKzcp
gqOoNC7yWXytqhLHelZ/mG6NiTdHqRNi41YwYPITMZEVe1y1eOOPBhmJg9YKb46mIWZdLIuibrE4
5qef8M4NtSeMeTv5UMxMDO9wMCqDGVyTq0YS1gOalc7pZYpPqEa4uWJwKztNrouogth4PdPzw0R7
syfOF7MwhAhvrtO8+ZFOeMNkcK7pD2vcOjQhJgYMrYxlM/KVKUwn3Z93zQ0K4Qt7z3YyRJplGACB
i3lIBqJ6fAS+ugj5TYOnVwZRKKx5aaNeB4mZH2TR1xm0EtcnYpWVHVukocZikrchjAkyJ40oyYc+
P91iFwAdqtsZ2Ciw0lR2tZna7ateGHLxuFdzhteMW7GxFT1MFvR+RFJvN5aGiYbvxtsZVdcsIqy5
qizCqqzoZdTpAddK0CSy6yvICNuGxL53IbB/3ypezlnJgDSAZgH3hLyOZ0o7IjCCH+PWmyhcAGTC
ZZY+2/HP1/Qul8YJDgJu9YmAEf3mFdQY/CWO75MKzNUX599BJk9HmaPBXWx+U6uTxK78ZqROR2/P
tPsJr1GM3v1gD4uflhrnVYIDEZWxaxcNPH5h9Vk9rKqwfdLRxMFAJ3F7xNeAhjUCC+5vB6J/iG3Q
HRBM//G5VKgQHX2q3kvXm53AoD1QEWelrneFqnMMxI25v1FFP36wWGxdJ+WhsIv+sOH5BHMCVCv1
DUJIf5fN+STvTjFUMG+hYbMqd9ptzk/OWqonXU4ScTLCbWNqAgKszZsPMwav3Soa+LTMtWbwpTmQ
Ln8xBfIXmkWLi6KPf6v1IA5LWzatMXn4beQSixHhlTgVjrjkLGaGR7hsSLolZNOfZVpHL5A0p8X1
GCX4IiP6O3nGOAa86z6NNpVDZ3n+dSm6Roy+lKJQLu1lVM2s6Xgxsrcb2tiBEL8k2i6M5xJkf/RI
JOnzNo/k5lFGoWsrxxFta/04flMhcWVceDCyN06iWE+Nwg2HuCvDDrf6qcvem/ttGvWiiaVIQcvx
3gwvC96ADMutPOsKDkFrHLtPEKCuZVcoKzcQwCgKdf60HDrACQlSlvNNasnm+qfkh1+EQStsBx+A
vbBIBK6oUmP1Fjqw+PyzitmQDYhAhvLBkpvIkM5mMMPl18XjXj2ZTp0iyVOtCFj5NtHHKjF0JbkM
fUtl3bQybBqBBP8uw4b7mG08pRbKopXZYbXcka0Yseka5uJ0MPT9BGgikAc3JvTyNDHKP6aPKOo2
LXDLD37itktQ4b6ObB54b3vuh0TwBtT8EiU3BznEtgJl0tz483FHNLRj/nY+JeXQP9ho1WlcWWof
ZDLmlve/O2uSUZskzgAJ+c5Yn2rHk/ESMojl1dbywYKn3uyLB3S1+dchNCQO3b4atby6k6IQkpIy
Nz4LiWPGT5P6xfgBoM+K3cvd3anygo5P35vdEcZAKqriOQxio8FMbie2ZFfCdd7L/vC7ue6Bwx6R
AYY/Db1stGXYQxUfQXVqeE96GNH7yJZ/IpFDlOC9rsDOYVcbpCNUWMTL1TaNMvRiotdYkdf8ZaCS
6+Qv7SJFCxCmNnmBzSsXh5JyeKG4O2YleE7hS1XZiLGvOy/rpVY6lc/4G8n1SCCF89k0jNk0m3Iy
wAIKsqc+EFxSkxZJ6j2hb8q8qYS71ml8JfUWoCYVIsxGv+Kfejgbh845XFqBQdVcIynTXaCVoXI3
IZZ8mxx4vDKDLzbwWrndYnD1YcWV4vD/QlLoaZKlFnC5zSHS6WB4MjaWLn5fXFE1ZuGxVFTfqflc
h6eqQjrag4YLIFdDKeRc9f1qTh9giGEOiZjeV8EwC7HTrgySOCKP5aHpWYxIcS9+0pWar0Whumqr
cHIb2+niQqX1mAhJ8Py3Cfb75EpULM4+1jWlpV6pe02ZR0mIjAfBIIl+28ZyXGGI8QnlKaNSXTxr
R3eBwZ6oUWp5JVpulCYtlRJNFcaqTQSHEWv/dvC4fmuHem/6+g3frybe/Ev//wtIbzs6VTS6TA1c
XcWvEqjveL6evpwuEKNRlDUlcs5ubF+Q9cngCaEhqjkpzb1SLyDw2SY9lFDsqZE+DAteYmHVShxp
1uCe8qjk+yd0baPCUgDMdXQUgcNroksSPjfH07qYVAQzik5R1Y8cJAaUr2KeQHOc0ojFclHqCyyb
1zA7duAxYi7OLoBQFxnJoSx7RuR0vza8Jo7lBAaB9vYwoLhcCJRtxLMUKbVdEwf2kBoqW3yFgcQe
sFvLvt/iE67wNOF6w/xDYWrqh8eyB0iYvdxkwctUjtl+fJr5P/Km7VgauZPXxRwxVXyM7SMRE1dD
kknOoBb4lmvhjLQWZ9dtQmdguvMcYidbdXeGKQpfryD65BErrTja1kmYRelDnb5yT/68ZSkw3zzH
Hn6wfpjBfgxd2FBORRRTBI3axcNeoClmiLEMi1U/mYEe+WKrQbwdpB+aeHvbHyGLZfJkm6DMVq5C
UYTbDEhO3OlpH7mxZFrxbcLCnoa4+n4X2azGT2gfD3y3fS1pu2VXUFZTFDadYL7yRvt3dOBlcYEz
xfQ1GxWQg919HITA4n6PsbHxCaHBTjqA3GbzUfq/sBmKbuC5iA/w/13MpCNGC6CioWRwTGHKA8rR
VhT0YPG6dD/6i23ZdLIja6AGIWxQRUu2impVEPjl1qlYA/XUARQBo4iiFFfLkfSkVpeMVI5nclB7
8ZpsW+07Ze6ii5QEdMNesWBUcqcOdU145RjVYMp4+Zz4LG9W+sNuZLpEEQFxE7f9k2RoPo54VoTB
9tj52y1zs5m3iQMkg2T3tVfPv5RHUAMmxeYgqiyzMU1cXRpJyVw+yzfy6wal61za8U+vchBJW8w0
KgiK4uBo/6fEeg0Gd0e+HFciwZIEn9dZs1ldsnxFmdgC1QBMt74KU/EGSpUMWkCWvSFnWw1LDxkI
SeAi6B8waXjVWK1hbgIjNLGdqkTncCSP5ExDB8YKzhgmPMKpJ261eMqnTY1aJQVLcyDaaH7bAxGv
vh0UcstNi4EawmWrArFCCVSD2njOIw8/SVW+FtqOe/mchW/5ihax7OSrlx/8I0qSkhxgMSPJCXY3
BYMtcAhz863LQ3CNZZzXfxuYTuVfHfT/HFhcI3A+QfDHcbb5NPBl+OhpM1beJMT6OgLoApbif3lI
AlfsjXwgIdaEa5o8Cb0kRujdgPjjGaolvY2MwB2oSCA6fEe1x2hvnUEzrvzcSN4RdFuESUxKSqSM
7St54lzK/8Cn1hjJADcT0KdFVKXg/UDl0eAdgrSroJa0baPzTaUFIg3pLQf3J2SPsGKnCjG3SY5M
WCRTSVB2CoKFBMlf/k5unpvxwzIed+R/CKb8TJ14To4s7tI+iHtliBp/LqZVVhSqnjKJ4ooj0Oi4
aRVm1kNnX6NswESVrT2P7qtOm5NnA2R7EtcNKa2/b0gpoMv1LFavr47LJ15ogeULcmtPpDTPZGp5
mvzOZEf0OJ4us6uLtUQpY4qSlNJx3W8f+24qZAQ8La9qUeMjWTGUHfuJeyFOOnQ38dfFZ6PR3Qy2
TWC0d08Gk0tmIa9r7E4mLWm+9L8AB15Rz6KUEIS5RkAX8XtRzyAXcotYa5jsKCy9lGWMDIoVxNH5
qD1qIrkJLznmgk9qNslqLPCJCpya5454CnWpd/BVlWNWdSiwc5MPORFb0fhQf8fBiZ1qfMlFTpTS
uf+lHYy6vtbfAqoHOaUPkU2Ry0+SVAnJxIu8XhIvuU/2Y3kKwJcorPxhnmRqauI2jRWRlAbIU3vX
S845UWWfctg8nMv4oWKQjxc6Ye22D9yEAvwKF9ZpGEjy7dVYy5nLB+wWX3UlQXoAkhYNLvdo2vgF
qlOLVlTuM7lVRbvIxpj00nJu5E6vT3mjLemyS1M8rXJAjgbISKW7qBgAcpbhMzdV8BF+EZUiWKTJ
EdDYWR2xz3D8kC8lIGgxdsBZV56pLyMMIwoT/irtKvY9IIhjcaZ1bqe7YEuHR/R8Ziaqi/UEuEsc
Em6ZcVHQqCsKmdO6wRI8+BhxKn/r7xGo3cKy3yqUOs4pKHhoxUkCYzqBWM/QA9yg6OArhfpsgMmb
iLYuob/ok+oxeKuZGD/jL2T9eYjMqtARmw+h/NrrHhyNdVGW9xZWRhYhQ8DwsrHTlGneMgYmg21d
OqdBa+uImXpk9B5zdwQcAgHC9A48G5fdDTE9LFNUp9xpk+VqUL8/pqIL34WVM0vaatMoxYRCr4AO
GnRzR/fubiALWOUKnEo0d6JoYEb5zuohzol4YWxD3voWXPZKx53IrUTIZ3m/aC8mP4TqzOFWd0Fe
icxhHzY46fYR5PXx1TE5o24QfdXzJGGXQEcGHNHBTcCsJsX4WK1vU4dvgYS2hiCC0f76QmMDaeoT
K9WbEwSyK7HnEDFu9Ea63CRF9mbhMXEnZpes3+WAg7K+gv6EALhudSKOZMyxLcnAmqrmh8QSG98J
l4n5A113TULz+1OtUZ5Tpldz87zpt3XhECCAi2DGFri2wegqaRuNAxlXz9gmfLs/OhbtIELT3LgM
mbXf9MWYJlpI3NDd1bdNr4S11T78sMTQfCG8eiR92IMiyNYXt3sy6k/OISXEihIBRSEfoJSbbJwQ
lvlT9H8UPoXB2uX1dZmS5R9tpiRVlHh8Mr+EUYlQT0JAGV7sm191iaWnBKX8O183ZOSLJDMkiWoY
k7V09Oao7nNcpGTpQ2SHdaOctSs/w2arBglm8TujmV/XoLeqrXF5Ppu7wymIHAWIRFFCymt4m5Tq
3K9vYBuna8QkqudXV7M+3Hpx+C3+w+3ckvg2IxrruaJcUSzZnXnQI1WieDn+6DksZtgRd9txqPMR
2ilGuD30T0fNSATQm2jYyMwKtCc3KE184UMoWto/aQXNt2NM1HvZmBYwoOJRBZ87Ez2d/zQIdhlb
5LaEUL8ibTBUmtAx+UhYxzB2nEBxfk731B1dd3llpDKpiynuB6PS06oibRE7VZLYOQt7EMM5L5vM
QmYRFvLNz0TvsMwfANOAs090iKl//NVcBAK6IbrH1wcptCHVAntXfJI5cU9rkTNo+RV4NLhS79yk
AsphWIRY/ptglM6ynXKjK8ejDt6F2fP3bOIgNIwqqrwfZxLwC+kAYGrbI6OtF6Eb8q+aAbr64oTN
5osqzTtTxLDs7J1HSgVPg8P1yHL7cZvUB9v+9mMXUbhDH4k+JziuklQPVX+7TL9+UstVurULBUPV
F6O9GWOJxiZP0Q8WVw4+Nj8tFokRWzeOz5+SdaBQ3l4r+Brh2HEgIH2HSqMEs2EDLoVmYEXa8VL+
WeLfqQHyxERVqUm53Rb3K5iOtG0YQsvayH/L+5LDsFDMxMHDnH1YJQwngnc/4Yz6ObLxHnEKya+b
vnzSbjyWPakp7BHpE3ubvvR5Vsj911esVU1Qr20UvhqohnlAqqfvrSCNSh/OTkFZuEx+/ql27WYw
gTwm+GB47HdtSHHl80o7NnnpkzEYI0HUZ//aSJpKWPufNMGn0VjqvLHgFdwtlnD1441IpS6/0kuD
mPRX1hDTQ2ia1WD9s7KYcc/OtMHZ7eFavSoafsEmLFjp0fnoD4Ri1xLV9M082WbtOWVaK2WGpPq3
gxe9pxZhzLyTnbI/NQ6lGebNfjoekMH5nVSTtIQ6LxCKWgaqyGCfosgV3ghbeXK4IerPToOzUy7v
92t7KfPHAFw2HLzTPLznf64enbUamMctUaIX/pgOhv1HwLmCnthtBHECN9V7P3pJz+VSV8mFb5Wv
LGfHiYnKfIUu90uGpxLWuJ5zzkSrM9TFJ1M59+i0C738M+Fy9D/ofU2ntza3mR1EGSAd+z6Q9cLy
7MBsRNJFCdHpMshLKK6NC85Ke1qO7XO525ryKtrk1+PN+g22lAIghxj9W5LQhduNeusOqhy9kY+U
geoK7EEMZt5y8QjkPG5ny20TFxgQ7q70Afv6k9xLsVcQeokCKiN7xrOuoedQipY5GT7bkHJCIbmS
Bvnvj3H6f9BDNq2gi8gNZ6uO0VrGkiYMPHj1AkUmAei6Jg2LQnxXnO1SWrXReZY6/+FwNr+NNblk
nI2DhterT6fdWawOfOr5q+rtOjCS5rZvJw/Lm9I4IEHQZTxskTdSlvY69ZG1SDCsTl9CF14pYCKi
IlWOoCHPE06mIC6DDaPvH+HfPfAJVxv+MWfphVyneJOiSC2uqzwHX9z3/5xbOwFM/qem3CFwMldM
RVe1xoP7v8E4e9TgrScxElzhVwbUVXF+hd4jIXpCmi87WxD33pyL+EeJl3UCpuj8yvAnnbBHqFU/
PEDTcwKQyr2kLUv3Rs45SXVKjRtoMBkuMhbZFDUsj7k8EuKMR0puoweNESs5wWz1q+cTSUEGG3f2
tSGozibXi9wP22K8Axk+PmLegPkItAJkeWFDL3Uo/wpEi9BpmuaadSg3hpLa9S/wzL20HsACdrF5
AXbxY8cb7J2T4CYypPNKDJ6P1bzpKYRnXo8wy304gEqFr0QsNJo96cK5UJdCvJKj3HHkLpZUY681
aN+hNglmgWjHPdmyluPRNC/Ip0zLaXwMujez0I0uIb0uLRw/qQNCLwnL4PvrGyfD/hPnqZFSoZ9b
b5SyZfN/BdsvctLXSckNIhyJHaabT9yM7O1aatNFwfRDu5nJeqZ5O1nhBzg5ePH5HAsI2o7pf7fe
27PxamrV3J737r9kQND72AuvZG50+SzZ9Q5uphTaQ9fleT5tMvKk4rOR4cNiOEl7nmFSEiRa+wyn
QYWHyxukuNA20D1ldPPEHPWhYlGuOdYia+gsKjYVlhQNsxZZr5pwxsM3sf5T2SzkK+Uz1klqQV8S
UDcAbkM6Sloh+7i8IOrZ0skMefbmXmPHItUi35mpMrHt/f0XoZA/71PTktYSYrc/VvJNLCmkHZpv
fWU6Ooqsxnar4e1PEDAIrRBQNwrh6lRo/txPtKtK0sUqJElQFlPmGdakHfK19TMytdbvlm4fqT2u
J+KvLqptWeRD1RZRH10ZVa67Fe1QZiUdDLBGYZ5LNl7KEk9yP49j4EGRn2CaSUkPNjav5CksEOju
v/28ymWl6Gkx54w8/zqxi+up+SWuczTNrHg0nyDp7w8aga6jQaAJpE5/ZAZ/OMlex37gpLXforHN
Jvo4JUF8BFHzM16MbaEvvAiA/rmZKmqMNVQIa8ebfb7pXkY4OptOOpr9IEecIjmZ5NSqt/yMs3e9
8EiASE2CBu/D+8Ty/cUz4qL9h22dktUnEkYBPArm14z1u0DHoeB6BGxxHxlfIbBwRpECVCWdlG8B
i5capuiKiGaivnQCx5CUjit53cJuUqnP+/OclX6EsqlqqFpRv2GgBTyIuwRlPtquCG8XWzjZeabZ
kM/RcS8CwCt6yUzSx4P9advYx3395JR2Jrr/GYyqSAsOumPAmvpdwI3aQxP7wbJTpe/rh3j4dzZd
Bxu9KxX5Mgue7AHqRzvgRXsgZgxVFM6FxCM7vPFOjrCGx+OmSNYnFl0mFLHfBH1aqMxK2IgM3VO9
ZJlqH+i1AdyP4wGkcbzjpr1lXGn2r4Ca4ZPZPpj9xgj6zFWJ9T7hY1KvzKhXrX6rhXnO0blbC2As
2Wehlai7Gc1+gKqSbFzUF+aRrZZHtASY9etTVBMSBPGi+SbuRLKcqYskO9YOVpEc0msqx8wi9a5G
XQrZp5RwKgEgeDB2tvO35GL09aFl/sp7frNpZChgrUUqwXwwx1LEq5GdtMYkKTd/iZd767UaUVW6
JtrCNYaoSFX9oqCufRQFlh7++W09F3QRU5H+kWKt3D9UhhKcFoLlL2MKKMIC4BaCXAwEXS71nPQB
2S9+i4omz2/cfDIiQ7VTMe82WzdCJeN4XmcDMYB4+RrFfh+K/WrwXCfTQgkGtmokuE1ZyHnwXSoS
RlrtUAPxWnHviv3kWfgmsxV+uyqnJ7CuWDdBwXo1VDfoKGtvKzY7EOpRrC2t8vi/zc48ObF9NuOx
U2rNXaX8/kum3QMwWZYe1Yhx9CptrjVPfdoJI+eaA51erOnxCG5xQbWBmTBzt5zkvtirtag6Z38k
HNg4cw7r5tIcKcZAKmnRsjhrrWQlHQN4le5ZbSUsy9pXRK/7X6Dey+RDPjLKGgDUCIDeQL3MdIeB
J+MbhNzBL9EF8//Urp6LjPV8jWk3suZSG4XGziuFMRFSjKUdeGJl0xj6rU132tAaI98pXHhdB4zf
unkv9mJxtDXg/EqcfWcVoxeZK1DrExmi6cELDndLDImyyxVjbLT3gXcspmR1FkYWDKWV6No+ExQQ
kSbN/rO/Ba+jZ25sXXZc+1MJF++SoGgkQTropSgFvYJzb2VA5xDmEiI83nq5iE/yJFViQiE6ISQ6
3CLNcM2XMZ/2IYEpMga2TXe7T9ybgNuiX3jOl+De3aJNN3qUarZdS8CEjxQHGEIkeXimQGdkenmw
/IUqhtmuL4qwFmhlIMTRiuARbCPH8kvzes0JckvjYoGmXHn/39b7RPKJp7PGI754gmdxNUqXDVfN
spanPqqi7Q38f/mTs/Il0Tnphab6+E9SZM+RhVSruE8JsZKkk3EipNXC9QNF1J5tTT0unv48VwGG
oUQqFAloXfwbfzcmAUEz1CO8xlcvUNPKEvLs4eIgPy5WhJVJibkYDmjeZWZux4r+aca4WOuAz/6y
xbmpz2aTl/Resb5wV8F/7f6gN84jnfeBYGKiANKmDUWDezNyyvHjwW+WY3DEUZYwgkJn0sRj3Vrp
fA9fKGsaX8SBNe6THU74pVaK05u3dOaaoYgdYERXZRQwOgOCAmdtE68APcrAS7umy70wWjCI/VM4
wn5CSzEboGppYBVcCi8ezPfuohbaryt2A+/xiqj2Ey1rXrZOzecu8RsT53ZTYs3Oyk65P62snHKh
iwryvFcOYxDuLnqJ/ELtphJfi5bOyzq3QvVTYyCm9TUdU9JtkH70KZddJXp6s96gIy+rXNIKYE79
UQDU0ZeWOtu/m+RzixSDLa4A5q4+C1lLGZIZ0DhH1b2FDobUrQRUk4P/HUrKSi3sLRsDfqi5S3Xo
JCqPr8ntELd/Z5HQQfdTzy4G2DGANpylPxGSSSLC9LCsa4K1Ki43pOIZyte0voQwy4ozgWUvx7Sc
AoGHvCm6jd+JhH2NqSp9bZ8dw7L/S0Iskldmh63d75NfH3AZXFl4xvkz7qdtMfRl6cuAGEUcIpNH
lyl1gpQY0vkCp/ufTiqcBqH/AXWREFC0njTItdOchb6b3M0sFnBrNGnIvzaNMRi5G7nZ273vJDOB
MJ3Fdezw0APIPEam7CYvFRZqqSFkqjmdQBolI0AF3e+g4VikgKuBlPBC44YhWbviP2vus/r34XDr
eF2+uHJrkGNaeyK29BIFECKjlvBzjgl+oMeM6/pWlNUZLTS7RIByK2pW9W8+QFJ9JFo2p8AAaEdY
Q7Yw5shmd79oUqteiFeSDmAuNU2GKGm+gauCfcPBc1K23FpOKn4dDH4brzHalsrcrVjiAL3D8CC0
di69yJ/uHpH23IBeCcVmPdsA76HHx0t//inIem/cz/deNXQ6Ebj5Xl6TDcI+jTg/E1j8Eiuo/wBe
KmgEm6WkzW92vEQ7Wm7jmxiNQ3ECwB43Zv3lDfYlFPSvccf4Txom5OvnchaLsQ1OjfJqJGYZRVnw
L2E19h18Foxz6LBN/8wm+p+lg8p0JIVl0OcehNXPvaMzNKyd5xGQWfJxi/8EQWVuP8QvZwxJT4Fp
f4idRBodCxbHjDPXdTkjps90+RfOefmrU7L2EnnP6FikeVG00cfqlnA68LvF2FIk3s/dJxeTrlN9
oe1zv60ANttWjf6jkeHNFcezzCRqk4FoUfS1MrzngB5M/kKDfXf4i5ceTqk31ymw13fiSvw44dMS
XmwY2k3drTl+YP7r2k46xPfC2fb7prI786P3vOJuyhhqjYubFsS69qQAD0FLZtZek9uZLQFwLYk/
KeXGUgIxsJggnkLFUxGcZUy3TkgFQ6rwwYT6J9FXjh6sOZg/+vlnlmKiSeaxC3mgHSSHnYufutBy
K4fgLP72zIu4bGKmsIXFD30VNmvtV5Dwc95qmJzxZ/dQ5Loo6PELsfNmhiSJCKzJO6T2rxye3I9P
418Vds6Iusu0ZXWBPt80eWA66G7Ot+CHiFIhdUcyBqAiA0bNEUD25nyue3X7jI8hC6PMsJzmc+ln
+vyapamJWtD1W8jbkSqhJSYxb4XQjY+aZByxUONc93b7zfcNxrjbd4wpEhyDToHt84mVgGOBOU+a
TmyQTaS7WyhGbnZYnWOYeI9lglvRGm339cNB+huwIln2N4rVcy8fiLtYiXbuF7gSs8YtXBsbCd5e
MCPoG7a2uTngaBpXQPc+5cUA0sZa7ns8kyFdfnV3bqxGTkJIQDX/OQ/0PXwoFdQjlOvG+UmFaLVr
mZUrU6JxJ/pF2R/f8mCH7TfEdQLUGlDTkdpkkN6g1IVxOOslXDHmww9wwx87hrFySFgB/Pll7/OU
vrsiUJJSLmMoYnz+IRqFhWBaE1fxJ1t+iOM8nx7CH06FlpzTs4j4bGz9NMsj1d6kUqxoWN4o+NRf
gk4l96PzrPMu3BK6sax5Vhj/7TYPVgJ7UWxRKrqJolQEQIb47nVxnXA9AdHURSrNdGXvXFcet04+
HJQ+EYgvyYKFUxGX5B+awnMXUWsI99ZJbkslcavc6sjHadK8+6hSGJyKw5p5UcsX2597tXdzEnPZ
u1QuP4+GjvqRRPLoEEgofEFl+EykocKxxcKtlcPdVl1/8BLtrdzp0ch5p952+JXx3vbSoMMCuO55
5G337f4UMI5rifWGkcZkO9s93RSaqHQ+SVNSKgmENmtMPDrXl7JqI1w6vCnbjGezanLNDUhL9CWZ
Ecl5mMzMnWpN8qxhVtBJco+kE/5p6HnPbXIoBZzq3VprHv/PBBQXddb0kGBeEYtEdVzBSw17ViRV
gnNU47pig/rLPcMEndnuR9gzF4JauodowshR1DxvgFYyhnXrIIooXJdbR+dbXoNCcN/U8aRVRP0f
7lCHHpim2yPER6IpBP+mvc7/HJITMTviHNF3/pskym+aM4wk2kkOGrIqiSA7cP8QNJneTsz0Xz5g
QyOWmcDOE0JU+pmeb6XcrL175uti/CTsKMaae/TDNdh9D61pfXVwbQYP90hlJX5lPrPbwe2hRL0x
Pvgyz4ws1EdMWF/uNN/6liBJs6wopS9JO+CUjcnx7mwT0qwni7bItb/TOmhlY4uYuchPPdRQUb04
aEG0pWwWt2ScInDljE0E+AZKPbqIzmxMjgVfpgcDtGLUYBKj3lO6IbM6d9T3pEzoIV5UEqHsL5FN
MyQd7Ej7Q3Uf0bimKv70RZesHzxgjNhIMgeNuVee9K4mSBPBSpmyalZbK+lFJJOysd6sVcfmYHxV
7hFoHThvQ3wWKrkhVxN28lR5tz0Len9Fhb4/Mq0GHGTP+L1SSBJaXYTilhJlayCtkS8W6k/U+KvS
LQmMVPWSDJETVy4qa9p5BcJ+BKRg08Q6eQ+DbBDPZ1dsDneorx5qvTA39W+kmoyilHsT1OUbCRTU
UY4c50VMVwKcxvg0eFuqsj8sWynUxqqkaHsdpkZnlvZY6nbzPTE51LMIjPKVHPnCUNjdL0uRyMX3
HdTUVBN7L4zlB7Fb621jGi8GFAjOM+rSyr3FPwtzsb2ReP8KV3cIq1u5KG++JbL/OkTTm1VMesIv
zQpiV53sr/GqtuEKddfuaknKYoMDkQFOnmUJx6nwkOTnkuRBCiV0436jmbcc6Mk4m+gyhv4Uqfj4
onjQhehbHtQNjPNBcmi7VLxP/sxUBnJrxI9ZOVHmTuhlCRe33yBcQquODXpA66G0GCcmaU3G7FL/
5eKtOJG+fsObljSemkCIpqSisZHxsSzcTftdPWSnsb8NnScNNUHmexy451fHmtcZRjCQUuZENirh
b09c71w8bb9BXDD2fKBH+mFsEAYqmGYLD91dnpzW4GWHutehhcHNKviDvvOiYKHI5yLdEPM2m4wv
+IvbPmt1GYuEViLo2uWdlln0WRkgZfsbWybVEybkRngdUetHVbC8UPVsVLhFFRQSebAQZIDwnfDE
XMnjcXv6ajvWf7l4rHZjDSDoKeE5dVZNQ+3D1K6AhKJ5eiS8+zcGIFPu/2VuqhQLM8R1l0Wk1S6w
2kgxuy83a6IjZMtSdx4LP453IaERMy3bHUTUD3LIqbHS5KWZh58kkt0Siamo2aa6wZuTz6w7Unzp
Rv6gHQoXw1scYATbGd54LVnk0h4AsDF+yPw2oXWrcyVcw0guWrCMniEnSVc1A9o0/yIHGMDXmm/u
/BzhiNctzCY97O2Ji1R5n4NlfaHjfN9hRk93iqWhwEKtGwRGDPM+GnF532tHLEgv3xWGGLpyX7xn
4B033XFvGpxUma85jp/oXqKsi4/24+SQ1iDwjacUlMXEksOM7ETwSBKPkChglkVe08Rguvhx2Vrn
mnDxAm7OupsP5qGJ/c345aZ6STqT41BxbJSD/Y20IcUrC0LRgCudlXS+tsFyGWWTUkbrtXOwYlHJ
WadkR5JnmgoeLzVzvqze/yFCWVawe+fYasrxMp6oCzMAywgnluFp60Pk2LJRkZzs1x3Pdzb8+eGS
pd6R7/o1YSLLUV5C54f5aadYBhPM1I0csM41kWy5uENtdiu2i1W/aG0sC9VHkvvowSgdmVdZc7vq
QVyYkZJYF1Sa5EdDvLuJ7qsxqOzf8AfBku6TfgSQYNyb15Ie3wErzcDa8+WaPG2DbWWTVRtybm1u
JhXupvUobfuTtjO0Iegj5stHfAPVIcQOGCtJId63+uSU3nQxglKMLqsSsf86UelhqUUJN7chhdlq
14vxBXc3YjQeJ5Hm4VpyYrPGgK+O3LjQ9+IQYCA6L/bPpov9AC+fepZCGTHNlhC2uM1tc+4rupL5
/TcndNTEyueivM7W1xjOrJH3zRhG96J9/k0SkvAuMu5DfdgdYPNJBQ5pSicspacyT3ElihqyYNYL
38RTA2YC6T7aBQ2cS3NXSgcj0E+ZUNxwC4+IxHcUvQ8Cph9cKlHk5d3+L8E67n81e703cI0eCGid
bulPnPGzJI9ly7P1Mk/25ojOFcOcfu96+/SzLK8Z5RlrL7ilypVGCSbUue33cSpL2FBylRrBloKv
inQyeEaebEL9RuozNYsBDXiAiEO/uFOD1sFHWxsk0oZUvjqP4bu94dyNHlDo0fvdelJwM6swLbbQ
rPJ+1NCyr3XDcT1o7cx8NsPPoKFcsN+oA0ZwGfI84/9v7rpK8ym7JYymKF3r9aRPVxpGC6EPi9Tj
ReceE6LcitB/PMIX4ivhBPjB2lwBBlBDR1udu775w4q52uPuQtSLMAvS6POzoqBl5vbPMRy+GE+u
N8tXYFyGiKW5ltQCBZFZ9LpqRYkhfN9dCMzpcUCbyK+LDRyyJdkoWc2i7ZOjh9IAsunLamp7MuTk
9vWgcH40cQTL8PpzuVtK6fE8AC4r2hYB+UGt3i2nMkyS3C4qLTpjDsocvPO+nBFh6xWnCQuhBHjg
VscMUp7jFSAxz2q7lv0KNEu8nMIsK/z7kwCAVgEADXoxCHZCSoCFp6cwmjqUhJ7htH96HtT5uius
E+LMnnpoeRmsjco+AdSfZu4W/xOg2uLGp8fQeFmRH35IgahxabSKF8zITP0/FaQB4JE5xrbpcMvy
qOEI8rnIC9yEVNZ2k7kU/PjoOWULnRADhej3MclIag7V/g7gw9gZ9NGBUZZhD1neNoGbfNhUvT5i
8XY7HszwOV68hLU5lxcNK0JDgTtD4zqocXCx/+qd20RUszhRUWHPqPHRjAw8gmzdBnvKK0H33ovV
j3ubz26sivf61zj0Qj5rzbZVj5s5QXHqVSWNlbnxHkzHbDIkyBd+QJtIADthr15ZKwje7ND2fcFh
tfS3RkNkG/USXbVq28Lh8KvO75M5Duco6uxtMySFo7yF/6IzPlZJLRVfgojAhBG0K37F2Y0y4G6m
EDhUl3jhJKg0unGJs+3JcnEg5XwFi+sWtMHRnKAIPbIezDrESrlToUNSzonUrjYn9YYmgxp8itCx
aIj52bVU31DzMFOvk4gfNG9BrXTUvMLAdSVBDboA6G3RWzgbYJ62HHZ/06fojWHdJGfMzEPABg7E
FULMQlwP/BdQn99Iz08xqIvZ1WAhqClNdoAwZzdCfAVnO8PiYud4ghJkkqFVC9hlDHgS8AZsd4vg
1vFB/Z2xHh3rTBBCXcJIYNfLGlKIqiPOA/aHsrXiZEPJSBcG5+maPZy1hgfbdCLL3qVVpXLfZROJ
aul8qUT9otUgyDnPhNTKbq1KC5aZ3ll5/dJ/8J3JwnV/niVNqJm8UVfn47nPESyTKHSuhFnUE4xr
wkTrW9oCWq+fM1q4fcgl3dsEaUjYY5+Rc1J0BZC6yWQ2seKFKWjA/mZQDPI0vsj6M1SlKetZrTgS
AHOEifGP8GAnxR/EhQW+xxaYI1c+CR52tBsyOYFUYUeW2II9+5IXFQe8q4PwsoOCXurZMtEz/NK1
KFM5tbBqUNEO4thpwTlsEfAyUYN6a9UF33VsukIkTluHKqVGXSCEbL/JHTLpKxk9nkF+EFLGLckS
ay/7qAAAqC5qmp/WzrgoVp6n0IPaT6sg/m6p71Tt5AMtN3bXTQXGMxWHK5DpKQhQ7JH6oM7M0SIw
gphmyM7K0tIydMsx7rZk5JXlLNw2pcEetbQIOTKRTWs6uTnTjbsEoucbq37brBVRoDrqjNT0xg0l
ot8DAZ1kvsRiri1/f/2YukDrQiCX3vC+NsUB/0aEa9ofV8gO341LR0q8FTdn6sOh8SiDBnMAe8Dv
vY0wzVsHnV+yiJzmmUmJmyvs5eLPuxMQKPcB2poPVMXlB0XBhv7+9/qdu0c9W2qPfxR9OMs0lmUB
OLlwbjYUmIOK7XgF7gHMdRnqrs/hrtTdvDji01WUPhFbjHfam1YRPmsyYTCFWwWnRndwf8u0ZKhl
JIETDzcvHIUB2nuvetncRHHtvgBcZiJ6AP29wPRT6JfzxGN19ynhxtcw4hE+dIBH9HwL+PyjqPxV
EBQQyLA3IUwdYLBA6GKytQkR2oGnkPPOmw6DuNd9FhthjLsIttmry0h4ptZuBHsd5HIdPAqxjBaC
CeeNZAcpduzzoSxPhTQEVS73jtdJa5yMrJLaldZ9bHYvcDdZAQwdpyQSijdhGbIohYENoQdAogB1
6+vvnMsIdI/jii7AYy8YonkNJn3FmgdMJT6tK+CLw5I/dP0XomxaL5cq3HskeKZHhikwI2v+YXx0
Y4OgskKiGids2qHNCiu8Y1jjXh6wfBm2tFhOKetFsZC4w9MJrpdrJ/ZfCuEUu6hyTuhY4IU96D9l
df4nOzlN2woWYZUSoouXpHyfJAQZ7Z3FSPxxmRSdejoPCTvknIz89ht/WjlZLHrV8lAqxtSeFHjA
n9SBcDemUlqMFOrpURMTfeuog9FNRp8oNFVOG9mhJA3U6ZkaPoqCC40e9aXThjJqK/rqFXzpE0Qk
c7z2so+c4OnnomBnHPuydmYnB3zYQ9zYsUyjOvhzF8QSZjwKQd4ZcPC3o1ojrkwQ5LnGV4+00aPu
WMISyfsGXqkl9AkVwX0rOeW+nimphTISBL658TqmkmTT1+ToKO75hCjmvoFRE9WU2E7Vp/+YnARR
c3JqVGpx+E8d1X19D5pqg3rz81p5xKLso4yx3VryFksSAEmL+tGIPtIn3lb4DzlSFOZrNloN0uzm
DcN/VkPgkbCVIIoU0xaeHY1StwgqPSyjR2DEs5l32FH6n2IYuENvJzUsmZxJEcNpPN6PyYG1GgdD
FDYdn6YOkfxxHzomHB+w98PYg2q7ahNVR2WOWtqfpF/2+F/4Rk7HuFrIqjJFACMmfUmHHZj9kCWk
cJcZjh03vX/YevL7ax+818u6nBRno10ZbzPtlsCQxdLPOhjBouGvQVrnAdy65Qr/cONUPkoQpLvK
/SQJ3tjRitO/P7pBT7Tkt1KwV0vLnWD2maF/uw24dPDzQ7jJP78qxj5YNS53ZZ8dCXPGqhKgWNa4
v69eq9ITpH0pJ364Ff2XSI8m+BFak8yv44ja3WUNBa4q9H3LtnP9Z9MnFOlZ9qexRE6M2S9zs8Mh
YC/ocyXn5ZGYYZPx9oJ2Y7xPJRbJU9f/+vX0GfisfeI0rc3hz7VFh3MxpBzKLfdJaIhpqz1QVg7k
c53E7yx5gYbBUGVT8a1o7+mI8fuB/oKMs+DXnFAdCOgWOkOwl5syuMHPFiy834jso19UFeFkWT3t
AIGiNeh8ZI9AyerV6bzLlBplcy0rMPMOcb9cze9H8RGV/Xpor+EiArk1dwIi07bhYiwX99HE+HyW
gVoAwPb1cebGVIRYubQ22oYu44ADKE5e2E/hKNkYt0o1BtZIlzhT0/9BCGDeDRYt3pUguNFl1CS4
dYII4Fra9mSFrU0hEDZWD3Jp7Kqnikpa8gxWIik2DhjGKqZQ8H37NbmaT9Ps7G5gKKT2Xdj34x3E
22KDY2oIsNT6XIJyRH+KG5KIC0Q9PM5ykX2EvJ35moiIKNg0AV4mcHivNPtu1fu9iCzvdCZpmbfm
r7/UN2wibUFzOIuky8LQy2H7jo7RCygdt0W0uKhNH+rsr07HxlJDQCJ9FEWp7dg9kfsp/Oq4+lqd
oWZcIBRs2Uz9v3omUJC7EgDC86GUoxiqKYwL/YhJKmKCHuJleGx0gtL2U7WeU4kjgsNDslmmyxqv
P3f4DLH/FiO4SpxK5ufwVCf0wWRYR8sf1lBzkk1dbOVSANlR6wMGrlMsuOfvm79LYmFjOeLm5IhJ
tzk581zV0I25M+nNcVhBDN3qeHga3mapoG9yORScxLQvkj4B/gwAPQUV7GToGA4XM3YQ0ONw05VX
pRUnwH0jJ6uNnZoBDqZH5q1R91FhJKjqmsoZIDI3mOB5AumGNbtJzl8QaN2Nved5lKFW/5TUrGbh
VzsRTW/LomET4MBcdi5r0t61znXBZy9OU7O2SkZeibnP/3G9sa7nTyQBc1Z/fWxLpLgrLbc3Pypt
Pcr2Pqkh+6UTmFzM/AIVMbMQO/wsY6+bdDv4WKUQK9K7sZx1OvsyNHMIelzGK5SqfnSaTh9gFH9b
eBrp/TODc13seUprqN4RZ2esFqdJySC0sH7SZ/rn0f/2s10IT+Z1OP7Tp5RuAWCEQHmvIblezhLy
Ttq9q+ShzNKGBi011U2d9zuNiUVMYAeNJGaTXyt7IOq+hynOuD2pXf3sbjXo28DhkE8fhXQOzN74
MljOlsPXuigC+eXtDGaKsXntCf9rqd9sn2UiQ+AOHLjEiEioakRexqux+jnoaW3JGjBJOYeL3+wf
gkVKTad2otTc3uImzPX/rtJyI7dkHJcIOdS99Yr+8zjzWoEPBVHmSy8GcOp3QAkpd1CjXX6bHSC6
3emgoqUQLByd/7pWASxd5OuaBTCuOM8ut+wXa+3H6GoNHd9s+TKFfjcB8R6czG8zQZylUZeYuRe1
wvpY4q8wIA5ZooOpwm8pdpo2tiE9++9nzn9spCe7dX5Q7lRTl/2oxdI/SvBnEN8cDQPazrKY2Op8
A4ZwbxXEnTgrn2iFVEdCBhzf5T2XJYhUwpnaQ3U11R7D+vxtcaA+dGHcfNMOy8mZ+X44gQhWqWqu
chnepP1UPzepaiBWll1p9D34Rx0KjWfUO0yajjmU0w/xhBldG1LNizkclzNbuipFp5hBskph1K13
AO2e/4hxAF/8C57wmbeKmoHk8X8gCYm6sYLJM9CPbAV6+4W9a9KB6Qi1npXlS1XL9srxGg/ME7lm
/mYGSoOFh42I4ZwQZr6JXNTa0KtPs2mZxQNvOr1Pmp4gohqUnFyf4NNvVe/+rTtdYPjTTAPnf9WQ
BbmxFNyLbbXsaNcVpRR6+E16Wb8JPz0W4bGnCtuqQ7vbv7lh9uj1MVJj1jdSgRoKRLRo1tMeYt78
wO2XpBVLEMZi71kbcPS5Q2PTtnOPfTIoel6HJeYABaUsa6rW7W2TNPWLPIKSm2J7F6aP+/+JfEy/
/asj+PU7Sqs3pONlOHeFkSpn3F5WY/+AE3A3o7It4UpXJDvHnC/J1LVhEYHuJ8j45d5mhwhhpsXe
qO0g2lTWIIRWgkDIrpBvbj7B+ZcZcMCjiuGPX6tF+zBaQGSdDbG98yP1ay4yQoY/UKTdCz/mF5i9
coLdloJiSZICb/qHEn0B+HsPYUORoEOC3yaHFWklq4Ghu8NvzI+fjs0DVdsDszjp/yYAlK+cdYYJ
frqjf2Wd2iz2ymI4SUiHqXUmm7ZabJi3eD9rkvTV2YfMRAUjjSpUOqy3Va2zRdI/czpTWRkKHBtP
p4m1+1wTmfk4I46s5Dk/uo8zmzTgNahxwApPSxNFePF7sum11yADUuZOzlChBSGX8B86Ry3bxDr+
U8AF6cG5Tn/3CpH4dnQqlOhHGxXHHGaK+XPX6SuXK2l4AkrxHa/TgkjaPsp6Hf7USPIoR9KqmqG8
NBhBWFw6Zq1CVh47Q4B5ignzWyE7QWeujjesZZ+GGOiONG3eKySYOyvrIO8OShxHLuO6ZLFtElYz
EzWXqiTAXD6gLAHR5nVD8c35QI6jDYaKz3C5Sb0KDMNTTG/CCFOj33FwnDER7FEy0UZV0JUA2l1j
CxH53LzvOWu5vkVwpg4KUIwoAp8TllyP4JoF2WilKm2sYUb3xVezwveo7OLzxhyiTLyXszjgP24f
SiqopruAeNDiNoprG6mii1mu5frSOebZ9EiHmdmw+VO8H9/YOG2e//eJdN/Hn9jubmZF78W5RAau
PRlwMMI4ijjQcc3n1Sd9dY0uIHp5j3MIjp7ljhWbOho9N7SgeSuoW4zFg0kWc5juUEr8qLEy735V
yEB0bcafO9Iwg05k9oErGJwL+W+alv9BLPCsolS8cxn0nhj/rT53iy2xZ0NnOalQ9JDafEFhWY+O
3dBooAk/WuPGlYy/63dE0r/Q8b/BBlm5cXDUXdMPkMw0jVIiHlftGcLpkLRmK+mfeFhF+hUzrdvf
xU/nea3qqCi4E+zt5ubDP56iBOS+sudL8QeSwCaE4BJT9KKa1oSN5w3NcjkjIdlroTRzZy+pBG2p
fjg6vNFJl57bhsuAjnS/I3YI/07GcsbyW561t1HFYDiSOdQuZSuHcO1Xdi4AQDn59OiFOpS40EZb
Kl2pgvXk0/xzsKaO9RHasBin6Lng2lIO3GuoVa2bcpHTIj+cCOtVdRviMUpujzLXR1/4IZhKMa8X
5X2aLoBq6pRPgEfOn1LwHhRr2dwI9QT5HSstWu8LHMpwRou5ww4THQ6baEs7WH7A0GkwSVEpkfgB
Jgr6Gg+CImsSt4yCjDp22nypvZ/JvtHE82cNv4dMaj+xFmU6lGOwd5ycOJm1q1Qv2cHWHPl9jORg
d1q/IuQgeBpjfUBx01yL/pBwgnL05btVk/TUyc3jg/o/sPkX3v0qJq4N/3+we7m1teNgljTQfmD4
+J9PDY7RCt72RL3GEQawAwdNHEfp3ADLh25OcB5m8VtIPcp6nX/9C1Fiw8Hrk/cpIshlK0IvHmBJ
YswcQRr+JA9BJ9pqLCCqNCSe794rtz/YJLYpSjaXnHBWJmt1QXq3Wr0ty4PpRybott/DZP3MX3o5
mcgY9VNRAdUsyOL59caJmH/rLNm4Kb8Xmo70ogwfNKN1k2fdNZmxVYHaiuLvxbEh5+todx1wkKNg
g0mDkAc2yPygXglaU+Fu4WTaFIwRjDpQTH4tBvS+TdXULafHj5YTFqqYYqK5stk+ePLCV4tG036/
4VER1afWNmClxmF3rZgo1xzouD5SFkDeYCDPyJubFgUwmGKwZu4mt96gz8I6M7VaP9kd9iX/21wN
yRUxXyGESawDNzq9x+klwPLZf++b36DKSlP19tMY7DFCNv6bjdFXWWLFPp7dpQpYLB7X98hHrTIa
SG4gsbWtipvLT/D/WZIPv1/ja6oqHcORWVePY7YtDUsWooSCuUJjqjeiJwh6edTSCdykQlBKNs+g
GgqRSO+1ZLOIXKRT32/uB+c9nq/QitOAh54LbSN5Suat8km6J4ZpNCeKW4Y9cVST8J73b/k7N+f5
gIZ9sd6s0Ie8IhA1Q5zlzl3D2dre1bKpYk/ZEadH1n272/9dCUvbGX6K2Vyip1Gq/MOIZn1iM4l1
O6KFDG52aW1GcIqIDhi7cz+d5GNjilp5Q26agPVSDfwxGORzHnQGfmg+itTlH2xxY0qqdEy05EFh
bapA5T7YnD9rYm5R+JYrviy8CRIkq81JR6ywH42L1cAVFTXFq3bKjz/ha20E1fVjrR66Ic++OMWJ
NquYReBCHsZUDAuoBPqpXdERam8pUZoAVBmFRegYUIcsHJPkijEPPbXKRZN7DyW+i6vCmw56lVHb
GGJo35srAV64b2WlbgRqJcP2JpxDPhfS/xx7t4bxzVU4rLQ+M72omcjGWTeDVpMoqkqgMo1/LbWI
gv06s4m0tD8QT91RLgN9ltSGGbk0KpMxVthhRq1l3gic2TCUU79Htcrjxlci28RjTqkpVSgNV1jR
fOR/V+C1hMRlnUwqDBsbddMv2s9EsmiaNdTDFCg+YQW/5Bh66KObxUmNh5n0cIzfzuSxcOkKbA3l
uCOBsN/wgIB8YT5wjYAChbYWdE63fokKrdoBev7aAw7u+Vc6ofmhl037cSKgJSR6KGi/hqfSLvlz
x8TOESlgoNxgeCWS73h+uX79AOcm5oRlHeIVlbdKOrlCqRBvvFKr8JOd+SkwDPtnCNGrIklxVxQh
bHZNGXcb2zlrTbbEdZRQcYUy0uo4dJn73XQtgiavXea3JoO5vT1dvYreFfl8o4SSYMG5dtPY6gYj
5By2uLJLLbuiUqCp2feg82ZJBk1l6zoXkIve+AFzzx/isnmo4KhVIp4BIfH3aDIHVJDVq0pERkuu
q0FEvMS3ySvkZu1gWhfOW9F773VAo+tL2t70Ke1bA76kOYN3f34dW9u7cCO+dhYGMUe0CUezRedR
WWYe4DU/4COkSl8LUIRtm+yeaCQZRjSObR+g0pZDo6UKBe18lCCW7ZXfgV7s3Pt7QpvfDaJYq1xL
7Ke36p7BoSzOvN8IAecQTCyFcEVPq+ELjb12UiTVgh5+70EyOsfpFHTfQEwP4bNXayAMDbqimsSN
lTWrvz1oMab139NqjJUzy/O1emQFia0z6/qDEoy0U2HQ6xA5R1L6hFlUU+kdCkXi7v51sPRpBM48
l7HgZBPCb5RcZxswNaX4ph3C6xvlv9UmO9Nf9C2Y0MNOmV5tb02yVA/Hc1A4winDxv/8MADnLAwE
CZ5JrG3kK7PrnBzDZOVpGkfBxItXsN8m6NzmNmqwgkZ56cvezQQ0mnMhXgvRrXTePUW2TWMi/89d
GWmxyGfvtXredzdo6SzIx4OMKCr8itQm7/sNe8z0tbuYloG16M7/a7SE+etffNmWsJB9t6vKwIH3
6osaeJ/CPvOBx9ZTDyW3sqzmz0KfjeYF8aENVRFPcC94ousSagMyFxcmqe4s0AcO5u4dqevrciVT
Pavo2KuPV4QcY35agcTlWKGFCpb7eTlkWpyr3YtkuLzzaaT5/UR5Z9CmspmHX+5G5FeM23zVr9UB
8RAPVbjfJ5N0X5OV5Cag04AiQKIx52UYjOb2qtlo+z10RJCP5Z/+RM58ymgfv6UyVYQa0Qg/Y7C1
UCV/URfx6Xck++7js6xUA9drEQTt2UQRY6CRTovc+mgOFjfwjTEF/CMECUFqiqIEa4Ex/T0LockU
hD3UymTrq26tHoUtlpUdaS66EiE47U3XAwzfqMD7Z0Xk+ROhzewaFoRVgU5GyKoJixqiHVuDqwoi
eo8F4vcB1Dk4yR3F5ClnaPzT01xzCcjP0QdUwzax/YovcPc2nBauq7QxYCZkVLoEZcYUv6fK4La0
VsFPCKNOxF/BP2THXpUvxTvOwHx0MFJ42I0kIqBPGbdnLf/1tGMTgXLwJV4zCnJkN1l5oQhP+U9S
FiI/bvENRsL/k2vHARHsTLQ4ycQ9UzCJq7V0Bek6IGJsgfWq8+x0xc93V2PzBdSI/v7t927CFC4J
fwNUQYvKrVgQD2UXA7wCwKQqOXzaX6miHR7a+jIo/hO7MQWrFmjgZwXYLu0VfOeJW71FxopuTy7L
ZEgy75d4HfiFwvelXRa7wHN1M65YX6miNKFxODhYO6lkbO8ECIWIoBBfFrqUh3bmkHso4OfpQu0N
7HaneDpnDnG6hQkEK1C1yVxNZxhjIuOXFLQHiIYHGvnaK51UAA6IP8qLUZ6y9//TRXlytsWCPxBX
m12n9tGd2Omne6HxYKMbgkmMdbxMNOJNhzo4Cq+GhQMoLejgdAnWWcn7BNzjy/GlH5p0DG+bNrzF
Ksjjw1i6PRByMrNjVgHYZ//u82NHdFnJ7gdt4kaaVt4QwdLICJZpoXZzsjKZLVrz0XUaD7foZksr
SK0VlP/iRqByJeQgo6uQp18JYiUY12lh3XbBJ9tHPt7NUxAbO+Ka8dlitfcIrHM3uZMO45vs8ZTj
V7Xn6Qq1OgGQKNzIlX0d7ypJpasPkHM7F68VszsP58BrwPlpTw68iGCuDF/iYRqHVJHICLwihSdw
iPAFbCZ8zma3htUygms6BeZ9zpijV/Wz3dxR1kPeDDYuIKE8/cJr7UiwxOa0iu7Jm+LOY/XXxpuc
ttah15nKf7T5KfnBHTc50ZUhdpFUP+8Bvn/rUUly3xzK3awFiqIyefAamoyRJuUrA6zkIEIm3v4a
quLFvlNpZtvWLzMCDhiz/GHDPI5BKYwpYfzYnoZYrFHLO6FpeWMQcdLf4DZ+jWROaBTZGNFeYXgD
XC69Ujadlzpz3vpbC8rg8hzEQ1wLRs7hNC4PvrfkVjfirFbjl0p2M15APukftA6UKKIjpDpuHUyZ
6sXBWJFXUZH1tBaV8UWBTENJkgkFgM4GANG7LM7N4OcSk3yWkSN2IEdBApm3nK/VJOoO/XrUQJk5
2ns2Awro8pNn1RE7dZbS4sgQk/DiHFTdFJmN2dVV9D/8LUDvRGLqsbCIF+0kg6zo4WnZ1z/Cy9kE
jcf8T4VWEtteVvAS30tGlJXKG7AgPQBF3HkB5rbGUveNP9WRRZbYJ+QWrNDZjxHSnBbiqmE0nSQ3
eRts6Edo/AFf4X3IGUrd2YBW7x6eYvo5l8ZdMyLQ9TC3+hTD+Zj93ByI+L7iXYQhCvAJmtegmaor
5vU+uW2u6iPN+zH5AQIbwhtRZ5JNm7J67AZ8E9q3nRzYYMtkykRvpa0UeQnWbM8LiedfW+yLsRyT
QmmyHA8aWaWVWnso6iS0oWCB+ICQzyOrhN8h6E50IxKWVu3HTmyQ9aGlDXs3A6NGHREg/2wfImQH
nqiOz2psgPaG/VHG3i1X3yXasiwF0rbtyZLArWNi0ou6QhRlWQSqjERlDokOSmaEVYi0obf8vwod
R8bgn3b/Rg3YJUA9avdJBKmViR9GQFneNk71sP04kVMr7ql8Q7KkL6YV+vU5zJIaJ7OfG3GL0hCH
DrctfWrhccz4JjTTZKLMzvyg7giHeUqAwXwwH6G/Rtpiip+13njF0pPPTr4nh+Gyu7kbGjrFwfrp
hQjpWU91eh/z5i7yFGqrMAk6awRpZUjEJRB9zlw66IG/CK4nB0tspCCCF/ZHj/1F29A6swIj4TAM
ncwg1iaHlkyCENMh8j1cg4UVA7R4RsnYk8mcf4FXIN552qFLhTS+X4J1xyWQduy5Qf3ksde9aD/0
+istkYyjH2ScnHTwFmQ4PeCJhz+SDy1qsFe/OOLBv4gu0m1uhNlqHfqtXB/QOca9DSTb6xkl/l1/
WIYflZOZdXuJMfI/wcejv4YGIemt9jSG+9iCKSMATCY3G7IGRIzSx7cvqdCY6WlU4f/DNQI3boDy
t8buax2kT5p+50bos19sibZ8h4odAEqvuSJWohSePa9PYRVI+8BB8pA2RckZWdMXe9qy70V7d2iC
RlcbpU4WsCuS6dw1qGF7mfSmMJXI4lFGdQzReUhSicQhRiqiCox1lfvyk+X4CtQKowZEkHWXYXK0
3PivJIoIoNFKKSgjgQe2FB9hgBVeaj8Jpq1dnwUyxVqvfo0PY5KUGJJR0iyzU+RYazcNVi3Pjssg
5rX+NpNucSoIaEowEUVh5wtaIu9CyBvE0VtRDzgcP5t026NLCEWjF9X8ERgutKQrSSUxXDB6WEfx
+B/LI19NG4NMt5GdkkOcW4ONeW7hqcLIiiZUQIRSQG35N8syYHUFUON1IbpwllPzf/ZA/E2SFJk3
OWQAUBhnfyTIhshpizWy+DqQNkHcFdPTIjKbk7CNcnCs1E1fNWKec3WpkSRJPA0DW8c7Rpjz2oz/
dXBFJENRlWuGK/2g9gSs388g54YakJzQvLJCMq4y4UHWbNUY11i6hAMigt/8tUaDR1SYOX+R4yia
mF6Rd4wmdYw2QoURtScrUnSSb1z3CvHUHJ3c6B/AR7QB/niRI+ceyfhay5Kelpgb2/zMvzMq4wHS
3hbRTdsjsAxRsKQaMIPgi64rC+Ln2fZME0q/LehkQy0hmYPaFpvmsXEEabgC3yitTyQ9ycMvGV8s
5PHvOZqRmlh7tj5xmAfst6qHENft6N3zwPiCO6ZqUnhSm8wYEq7zOrLY8fACk2eBrJ/3mawlChbl
OOiOv2US+UxndNMOKQ2gJsRQOe147UrkpclcWUxyEwobrKsbTofSo6q/7A88n6hgNKipTlnjdNCp
fwU4uknhStPVI8TK998K1YhPju3mvOROp4OxxRR6bHvoW3nL/62aay8dvQH9ZYhRPAmbTOexZqk6
n/ldgK1gdr9DRsV4MIRBULs9y1SD9bwuc+dBfjtxavUmk7u1yIu0VbJx5Lvpyf7y3mBpJ3hn9R73
4d/XOO9uUR+HAC0hlW3HqT9bj9fCD4RT716/KgbEXqjajfRFch84NdsvkYyCoNakMbmuO1u508zc
o1c1DeWqPpKT3ldRSb2dStxP70YXFk3180C+QuxlE6/9gvCQ74meG3IemMLto4XXO6xNja9WNMk7
2fp40ZlOwtLxDJOho+Uj5JTh26YQzDg1CB6YWWIxekndSsNEwlvLI+Xl05/XeDVFRWQTfgqVmnBu
G1MH1lxgM4s7tHEg5+qGeKRhd067oF5TdSiu9syyl8uYhWFembBA1NcKqMdHnIv60xCJuXyZmPV2
ieQuDEtS368GASdckQBJRKnZD0OQdMuS2X5HNkM+a/L2TejCBkXr/kkXmLiJG96B2t25/ZrX1aDE
TnYloCn4pd8IfoKLAsWVko63Wc4Welfyz+EDA1767fm2ABGJiWdMHqzYzEWggDDZXApAgc66NFSI
DkyUBoQ4BqF3nmwzSPfkMw/xQqKSBavdIq3SwcwPyIdzFcvpIwbMKq91hmp61/95unSz5qqomENl
rUmZDNgJe3CGlTVF7AmR26JB0Kqcjos77ST/2vL9vya/Zpuc3JeQQ9r7rGLp2aei+vBMZ5Mhv8Or
6LJxdI2M9QiQ1Gusw/8f3vibxz83S378hl2PEauWqYu9cMjOHX6WEUocBOfUBzRFkQPfTDma4/zw
qhJCve3b+awqJavSbri22cuEXu3csgZe0D02AshY9msbPhD9M4vm1g/BKVhUiwjssqeNoR1TRLP9
MGgcfO6VK0XYvJdAqr58TXJXQbVCvOFQJQrQCeYes9CwkgS05MRg4fktJP9/F9PYNaxmg3p31brf
jKjD7ZY4NvF66x9gjiyWi4m0fvD8vk+DymjYde0DRCcuibXgau9fn/x/124E8Bmw/Fkfr3//3stY
qW9jVP/3sQJWyrzO1iE4CZGXjXIh2XMzB9EIBRhj0F7ZQxFlBOZfIZX7ieRSe6qLywt6ekoS97lz
KJ1lNgqBVOwrLMz/txyie0iCjjmE96TOOV0C2dX24AQOiqa1b76As+aK9lI0rpY/1AAbthgsc6el
bwqhc/hg7vzzI0nbcqqVgUIYKisOVyiqcV2Rid17Mk3sOjyit+XW38L356BDd2zbRlFi3iyMF+ws
fLtjCIS9Lxe0jDN0tz1444M+7z6z6jn23fiVo3hm+YC9jbwYL4xdtGocuab9LUJDc1siYOrFhELF
z1QX0p6f1KoFm0cbcgS6JfAmUP95PBys9opNCiqNBVgKK5MBLPPyYN3ojfsko9S8zRyzPJaCvScJ
66CSHvIL5hAXUaQAPc7I/DjofPhEYBCURXPmdBKOVzhb3ldcD+PylmErg/kTGZwty3me50P9VSNj
bC5TfXZHFwbF/8VdrMFWAj9jPyVfynKUZTFCn0VP76ED7DsyPQE5ThLRo25KBY5qxCpVLHD/nQoz
G8mEqRBTB9Z++2Pnc88+Xn//qRJEMblXWBk4q94+5sFzkoRQ0guud2smrFY32PMMf8ikPbL4JnrS
Ivhy9SI1GY5EjsIBG9Ytd7q+gr1D5yMf4EFFmbZd/GB5vUJqcBoLu1LMIC5hNC8fE3WJBq/AVp+A
uXbuuCli6a++vtfHtszNZYNviMPA7K31Mcy99NShb8AOO2QeXAzm7dQzMIASPEl1p3Hqe+kIOcFR
8tmp4vEO337ZuwJj/3+OdOoE/a4cY3FkuNUo3OKAfRfWUxSRP9PXTv+KDMWvJLZChfwhHJYPIVg3
iox9vPuuEm9VJPK2bjhL3krKfVu+7lRwJQYnlc2AA4YuLq6itiu4+4aF5xDrIU/I2E5RRJR7hTiF
3kwSMOugeCzSIxtXclsA2drZkduOHiNhjM7d84Q+JDltUNySK565QnbbJMMvMyx8/qVKBgtaleHv
7JI5z3BH9UsHf7DL8ex5r4jwPXJVr8w1x1DHiONWZdkjUnBlrpKmIYJMRj0FWUdtE5hXATsUGkZw
c0DYuYXiGeLpSRdbE+NQcFybQ2lJd9I0fR0w942wT6z/rXqynVeIGQ8kNKT4pRHuBH0yiFucuslE
A3f07GOqJHm7/E7YEpkDNLqW5Vn9IFNa9U6aeI84Gp3HgrjBvrIebzUJpN1o1QnwR7e85uos/4Q9
DH56KhFJM7yYoyzC/bbpv+ij4K1wxHalPw+IU67fl5DtR74kjFnMS1kzSH4cSrrG6D+zbxo7uQvP
Ol2UF4wHH5O8IGDjFgcF5L+yaipeboP/39K8Xop4vcnwCILnLJ9R/1avL7G9GQLmJCVZBWivYF9s
T6WKEcOC4yH2UK8qz7nCPK/5rwAQCmijJNJv9Jf3TQyO3H3F7jlLAEX3m5b4/AhEZ89peQzdLDcq
iMJ8qFQtZMwXQBU7wdfHqYc5/CnkYucgBvZ8SVNcJvGXiouS1cK4UvVGeXXmdQiXzHqZKih7S/fy
8ICYGsvoPrWfrn92rZIVZbjBOY1H/2wghNO66EU1p4GoKnzWB6j4YsluqhFNexWEaz27NPk85xrj
aSTpHG8zvZ+alE/RAasfx4tNKJhK2fAzow7AK6z/o4dgWZLmlgz2Er0bZdmTrh75ImBfay+JRbSL
gHVagrk5OE8fYZJF2ghefx77k7wDwL9i0FYQvaG4wlh4N23Yvc1/fKc/LE1VVmGGHOTTHU156uy5
1xL2XStHmlNJFK/HvEIv40FAKJ2+eLn+6l0Mntg8gWDXB7BUV7dQkvopUFmB+v7FXSYcn9DNDECN
2bVskdb+IMIugCO8WRppdenYD4HCJjvdXOJoUr9pXYhUEOdR0OQIHmPmFpGnbNaAsLWhQwE2ygXX
Pw9RrgIJAVX/+25K+QxUlYuEwUJiK6oov7ak7Hb8YIeXk8ssv+v8/plLkbgQX0xPVD2Ze4T75l/L
CP+njWOqkovNvRQDYVdFCcP75yTSnzBreH+Q3n0RC+Rr7X0qBejZZafWU+/kAR989mIUGcYs/WN+
SkOcJO3matd3xswNECunggsWet8fHea+Gbh4mFhOfiV3Ls81wdBjLsB54O3Gtu9/yKXu4GxfACPF
jkUXE7o4E7KtIde+q7bJkZFUh/+acUaGPIGGSrLPvxrh32UKkqHNXm6D/RRWPjz5pnY+UZMJRdbj
Jw6cjRvKjRJGsILe2h0FC2ZHlkrcxpdjiqYgzxgLSRfXpBaAWPW5Ue1aX4xN/oq8Wpfkd4Rnnkor
2FBkDjT4p6HrEkT0knssTySCQJua02q1PDQ+wTASsmlPg/dmFLemQsM1+0RsDtDOGiPUEyr6F6WV
fYUhmovjfoRAxwZFaOsim/5+QKGbveHJUvbGug16dnge0du+jftsv0bq5DLnGJGJLLBrF8pOSPgL
O/aV0cwWG14N7EiywUu+LZACsm4gp2hwI1M3AUrA71ygzAEuL3vmiXRT1DoigzKH492uNwOMWUHn
ySAqXa6xKw7fYSYncDwZSHAvlrljoG67IISUUSlObylOgURV5aQx/MzIm3Kn6HdSa4Pq4M8cS/qT
i87rDIyEAD/LIXrPd5yzqGlVRin1gE28O0d8metIyYx4bbgC7dsenUm1EpSJ07tPTBOSEpfG04Tg
fbbsQOJDaU0P6mFITY2XZL87lxql6+JRANjPyNzlxvP3kEwcMk8JLtmSYAc66eR5Dp2p3GlIw2FR
nMGb3LaMkg3MjWDYB+oly5sHwyMbtkAB9/e7+Grs+IPR7dmBN3+47sxM4sPCAdPc26m+DF3CvZNu
XKA4mZjh1HzoToQdY1b4i/zOlfhH1+Ao8gg6OfDpZWvOMVKwA/jMgJxnCh9V92zzrWrb3p6iku6w
xVVWzAYwZPkSE25uvmMu2GUoQ3aMy3gpfq1l6/hv00dWKj95M23zxVFNWtMjfgJGnf/DWCJAum+C
pA3liMJuDpSNUvzH7cWca62dTfGRf+QoceMHSu0ij38wg/VwU7bpGQtjuOd0EZWxdluWwKoiz2V0
2SWSSacQAkXRd63qXtg2wROL+up6jetDxdNidDwH3Qh9Kf6MJTao+Qg4+FhBzAqH5svO/RsNS5Ci
TayOPNoNwlHtYoM4/ZU+d5bRLxsgppy6p6T5/6J9WMgHbo1ykXSulla40AnhkzpHm7CpbXB8J+CH
BioyvgSxYtI6evHStVIfN6Q7leE/O7PH0k7El7QKUR0bCVdlmCpPpCKcp3GINlSDxTJIGfcpiG29
UA3UYzmKeRzo85PwZptFAbRFIlwqkMJwmcjzZ7NV4clFTUjA07O0btH0sxftyDm8FpFW0D/6T+rQ
PUCoiql/Jq51Y6JAgOGcy8dbApggxDztIEdArJuw5oG5ySqkg3UK71hOYVQud0y6ugjpRiEZaGv5
A4JtkJ/sZPJ3gFFCyJOol2kpsQSs+w7c0rWpaAB0z7OUecbCkVvShFhAlgniqSSIHeEVWKhHLyth
gG2tW6z0tD/zHR2SiH0RndefS7vH3d+9Nk8rKmiAFjOXpfsoo1HN+yd6rBzJAftN47lbQVjq+7fi
v66p2tE22ij4g46tVkFWomViJZ1zHpaIjNsz2Sn0Sf9dBaQn8vAoECKiLFHaKiBN6ck8aIzarlDt
Mh3acO01gboqgzRC2ciJM1OISnOmEOD5KsbJAR7iC2k/rWPaqC2wcfHkhyPIHsFaNgblAhWuGvn0
CG7XqqPoun1rkcImGFMfB9KwriIN9yXkuf8xrr/yMAxouH7NZBD9hPEkg+AfWuA7IKyMVCUlJ5oK
1fXfWr1mM4CsIkyI02KLXRyJZqAZ4JNkHnrEStEwQDNUdzwOZntxf1yqpyZCPqzWSRvVsq7O3bv/
Tcdzyg5Ow1IGIoGXqCh7Jd1ch0+FOSneGeOTF0r/jyTOxa5EeRFkzpcBeYs7sZpKmn8tn4jCk4yy
U3gxnghZ2Ci75GCTvC6FCkhwS8Y1fL71K2Bjl8K90mxojI1n92BPBXtfN6Cv2M3N3lNHIKe3BbbL
PlgJTqD80PEpDtB/fgJjg3dKwPgzo2OUCPbwgssfvof72qmqq4kQehZNI1B20uaYMKkNrsOE5bgv
uT4PoqA27dVY/1YGUOzLCUR2GlInt+2pVd1048AadE1EKRZ56h/fUz2cpKv7AE04EHCRXqW4quqO
CoUdD3Mtnq1I1w3fl75JiZM+opIpwIS5/jFN0sk/4mnr/gd9aR1HnJVizucM4vz3C7oAEzLrIFoH
wRODl7L3+PODZclcmENVBblKyPorkUYDw2iMihQg7m4XymHj1jeJ0QWHramwSTVOwu25t+Aix8mE
/MIwGDJM6xnKOOIMX2nHcisZRazzpMCDVxRVt1UDqkIOSCeBnK4kL52pBBcJl0tVGJH/KNmr5iiB
9nLEPt/HqBTrI9z3BUWaBTJIoS3T/DeW21K960SHACpfJMyjgwqr+qgMMRs3/YbHzRsm0uNwGF3L
G2ZRCrSmzW1vEz5+eSYu6ZIHe+IjcRo8xtprX4vrvpGLAf53OtNWsDjbcMJv5CA5eEdG52ConOh1
LF+0dDtjmj8RNv3CnqtgvOuLnMOJog0O6xPjzirsucHDUI7KAmFzInrJBxbF6AVa8gjOodhsPfWT
Ze7QRtlLAvwup86hUfHEE7rvb/1VFf20mNiyIsSvan8tpvwHA+jZ0ufFyaHwi4StVECUVxxPpjac
9VCCEs2VR4u07bT9eGN/P48A3pAEbK3ylJzcMQZlByZQPn4kGZr+PRRTUl/DG6Fs2xapfF3nJOuH
rvOMhPojw3VhDYYJbAbJosafRV4eODjlmpgIkPx7EoFt1ajvc0AKxHMqvq1nrPjex+az1xCdsmbV
KbKskR7fEQJbPtFuO1q8aHTcqxDRbkpWX2PDwAOxG9lQop73tM6xtWw04SkeTb8UD9NYIN3gw1tY
e+p5yr/wwyGyF8EpA7372uObSnIJJ049Q2339zkNXaNYMlIDHkXQI3OxXxrB9O8URufb+0mhGLJZ
yC/DDEHfdPF6+2AVNeAPGwz0v7ugtk0IQ01DkMrcvhGty13mwnyQ6CGOwQbw4ifbB5giH6/a2uF2
D45LY1jAgpzjhaXpDK/eHVKHFFv4e0vE48aelBUGB7tKDJ6KWGsG0i58SPSulplN+uFETGyD1dws
SAo+rpYsckyVspHQ0E90k+Xi0Gns4RVJQUzo+CGPw3vPhMQL0p+bbUpYrsCPObCWPrgBsArrzd2a
tVLSSi5FaC0t/TrQkyxGNADIl56Oxa4vACaHOKbxmkT4vt2SwRh8JlKtKK+e/mniOc01tcVKVRnB
/KS/DFiuOUOq4DyeMgpgA9n17ozpOJfpHfNRo2+u+4NWmfNwhDSSB49NYmbpNNvENlC6PBxWTIU9
BWv9suuf4DYJBTQFe6747hkAx8W5njqnBzv8SF6drKZ+zNLkUTbnXyjjaLQfWj+rWBW9pNp2s6AQ
5Ce137ayweklrHZpJqMDXkLdJSTb2pFoIiyJuRtkrZS1qSRbxB7ks3LN7VtJlj+O/+NajC2wnRF1
pk7DGNtfQs6Ybtq9jygOAIE8SX7B67/DpfN9+vE7hJLdr4v5lr6uKdbCuA+XYKF4UkoegFILoBur
uxPmP4Wc5hd2qlqRFsBGcZcT9Kig4Owokxze3OWKpfQH5JKetHcjQfRtn73L4vVjluDXzGCIlLrV
PlwGbVWYYfzKLOgmpnzAB6cMj6c0bZE1F6M5qdYBbVsGf2xhtubH9MTO6q8T9ke9zo4lUuf0gkIS
sXVubARAbjX/tRvk8w4yav8Btxpwaj4hg5kr3/UgEPdD8kL+KjxN3okt3E4hp/ewQBFk6H/SwMtv
dwudJbt94kHaxww7XbXR9hXfTwUB/m0dXVKmvDgQ2KebB4C+Uj0G594VGEekl8vj7bKxiir4h4vZ
OuwgUXJfRjvQsbMZjj+6gSJphOxqfOAJ+gHpWs3hSE3domo8NUlE7T//RndMuxjXUMo9PWQtojW4
UixNyr/VXf1Ruvhhgb1NbQ6O4rbukoSjY/oyPmuZFo0NeRKJMdQbf9Wxy2kaHV+FaT12Cie5Oybq
VUa7Wjic41mdSvKg182gT8nH5WDVXJ7es0ovplEsuhWBva0fMoMWCrjNjS+23XqvN7/WLZ4fjVrY
/f4DXE2/nQL5UqTvbTEUXdMPjtoN5dl4c79ZHJQ1s4pZBdEtl6WLTOuEZPbrqhJjkV7tt4NAW/Lp
rXQK5AEC2n0a1JAmqehoUQ9whmrmgszCkxPWcbK6HjdAvhvOiwf/U4YB1nA7yTCjDHj6YHOO4712
I7MRHKwS5LQqkYjMSbAgUGAabffmynniAE3rkyhteRolGWPD0X6bf+Xj5bsma6N7ByaX0KnFnUcS
d2iQX5R1Ovo9UKIHx0JJ0sEOErTUpuwPg/RFRttx5BAJdDsZAyjOyu8wBiJFR7rBwL9uovI+hlF2
2leuH9xW6NmMN7AG5r10ZE4afh/v9ycG/eKjQCQwkxPVL2SJk9OcDfQqzSyIdn0iMTLmHtp0Ickt
3BONGJRaNZXOvBUhJJnR8dNbK7t3QwTYmUofSrhsbCFw0x9/vNrfad3Eo+LFcpssFwR905unzf0w
cQoyuNgT8STvjsvr9MGECsktv8MwE71/q56q6CVCUyIxkMJj6qfzX0OeHB6xkOGGM9I8HdNsi3qV
iDNLOtBlTx3WAPQkZni8PZe4hV8WyH0cgKvRTldkSyuIfuw7h86bRIw9m5+iUKyA9UmfmhcR2tS7
33a1ULEhVD9GT20Vp0vWVC4vs8dmccePbjDNZhc5fbnXfuR20L7pch7tcyj3QG9ralE7TbMK0h2s
YWRXntHe8dC9dSRV2QZrQ9yucMSQ3gfg90t6K0H1bIRZ0SMIS+f3C4HhiyVoLpk+HxkcwnIp5dkU
dhB5FCC516iLtM5HV1x2//KBH5+2CUr7JJCQDLV9OfYVKKAGV13Yoz9ra0n03E1VzkdOyTRmhe8E
RypyqDuitXSMnUj7MQolvT5ALjhib1XwscM3hyGjNSsQPx3Sq5rfhcggHXtHA9zfLraiOhE+LBah
bqKejwWS2VquKHDTdPCFq4aUnWAKI/LHKm7xbVCqfqqoe8dxk7kjzUBx+UFQIZgW50iglI/cC691
Sc0D3DtKssegc7zGXimkiUN8mwHqjjmWNZXygfNBUAXKb8q3aD5J5NkWwFg5pc6rvbHRz4UN7c2+
+dnjvwAJ5IlxqjaQS70L3PgqnVIr5rsqAnkuz5utVRjzZlqlEmATYezsts/ohSRyB/dRxXijWuCZ
FS7IzVvf35RsO6/Ck6KwivB5gt89zEPDiFpkVmXtMVU/Q8E4OgYxTd+i2iTjhkDFWFO1g13kiBx/
ltjCAJccIUYnHEqUtb9JZNGaLUBTQjNoNH9z8V2QhOT61qbLMFlW1gKHmYDJ6xZNzClNHXSuNHfz
/F/Mt5kCIq40ZBUDQsz40cW9+IbOw63C7dc5byjxx82XvofzWDYH0qNiYn5QzIphgr/VMnF2waOF
LgPSxGetNEFxQptBPo5DSki9hbdP6ENemu/0AU/9JJw17nEOiTpZ79t5nIzBXAL3glcjl5a5wIMm
ULonbH2t3Tln2eqkV0eHeFf+qpOdbIeYTWlLjCblOpOhbwB/984WRXNL1hm5R7JZHB8xN5L0N6TG
dMyA0yWyBLhR+2+ZDKTbbtg6ns0thoM6aRAtQrtpfUNKL+UDhKsdWTZ7Z5sm2Y79QCYk0I2xR/A1
kPVX+cusvExtB5p1waIP/PxlpXehlUEaRjHKcD9Iaz/EY4Sf8uLK2Op/lN7gyIbD5weVFK9hYrJa
Iuak+kbC97fqynv0T1rVQRB8WRlizwVLyFfTsZyS+ErrbDBPJKO2dVjOavdFqscqbmZruPHfKTNf
02h8VFJSQx8tT81i2qtB3+dxWIasyyK3t5UBvyha7VsT+37/6904mPgeO2g8V03KTjvVvc1Osk/h
qQldim0+rs+thxl9h2IOAL0aj8tdBDa1DgYw8e5HMlV+nYd7TELVzTCEAPEk3Vjlvsoy8pqFPbAU
a+vRejeX/WDfuYLPivL2slDMlHsx6ltFr/cAYVGk2aXydPCAbgY38rNwHPbWK6J3QoxtqxGpCwJJ
gRHAbef44ssgNBsfS4+5QBKYLKMKBimwJP4NERAXOaVTIEmPMM5/wmoA33EAnmrVrjHckreuFvFM
JhcIwE/ehntKDBeTCW5tgXpValRdWVrr8+0sehPtCbpFNlRTY//Vc2UnrUluYSDMhq7a/kFXOmLY
bL955UgwUzbwMAS+w8sO04NhSEQI6LPr52Ssys/fI/GQCN9V8+GJc5hxPb6DM1zEw0/UbEhRdPlb
snC/TRyqCMyZsxyQcGpnykEQROdy0skXwLnFAYovpH713qhbctOlKN3ETm+w6K7nKV5hntckYR9g
vrTGksCDBRZHYKnu0vtjvAAkLgehUhQYcGnUWG+nVofsnxcZnmL8SIeGJkaiFIMT75FmKVOuw/8J
HNRxfyJ+aCC5adB4SbvJLqin65w5N8X6fVhILfqZu/IBeSZb8ys9dnNF4h1m5ynbv3Hn/OqtmlqX
RWnrFnp898GowLpAPE6KFeAIQyGecJXrBqzZiNE2JM3n31QDAKVprjbRaBH4a3HeQJtF1fa2juw5
oGSyJCg4V+XW0TufBOwRjAj/qaVQSOGZHKJh4A97jpnjjoyNsskSSt3R9m/aP19L4sOK6/5JO4nb
T7R4zg58NbErGV9qmjlaaoxUJSvFFIF/uB2Y6H/wjLAtv7uYiwm32/etK6Ckbikp8SfUdkhnqATo
cIWMLXfajcyGis7V3Psc8seqSrqQJR0O8oFkuEw/k9Br65NtrD0SUR+/26mBEP/R0NclIA1WpSFC
Ez6hMxnz/HcwwQ0kcNG7YoEmMKx06rObjyuN1QPnpg3YHVvxfBbhYpCX7zJhRlcOTPw+zD2OpOKj
1yGfqnk6c8onSMg7k+TRFeWnFOPCbZRd25KuG+huZ3uSMaknUcJJsOhgCTi+He1PFkfBy4pyjRKd
l87N1GAmbk2wkvNZQJoyuvZUaHnvskfxquT3EdjNz3GFtWLW3KiPe7rkLPWM8Qz405npEi1iBjqy
QrTgQjVjcaA9F4M+PMNOCEHigP9v1nfJtZYXqxjW2mZVHh+6N6FL8BqIok2O1gXvIKbfjk3F2wM8
eQAxXncS9pp+gOCzZyzv4RsP4nPg8tzdohq18Nnwkz+fNdLFacQAjxwft4fwkCxZGA6aax679K88
0tiurdeKeoVX2+8EoEE2RU0rV6G0HEwI5XRV3LX9G3+9HIInJ5l+T35yu3oYVDKFLDNubhDkBMfk
EA1jphFpEZ5w1CCTm2bwxyFKl7ru2EhzbAyjVdZkBGO5kZvxM3iMHq3NPsztpiNW5Lr71PubIVuT
5kYXEzSG3bvuk0Sd3Obb2uTobI2mhszDeSZ+cVvsb9CaPLkGf4ZWbmgOvbbwcM1Xkj9rXjrKDQbm
WzWndP8HI/efUgyawJVc00BA8mAD8FoQi9FpWXoC49N1aQYFTCPoRxbZUcF01Pyj4bhBQdUfYwGK
5khk3WH3TfsaWryMi6bpJMub2ST9cLqlzDo5dtOyQ6G4fcYmJXrAZcWtF52y4LPIX015LYJjScsW
5JdugiTmhnOL/DwomsFOnqibXxhmDWNFsEDQyAe6tbkH+ARAMFH3CE+Bcls6cepi+WFpBsBOPH+L
nbrcHia0LuN/cwTKj8zex77oAULdg0iwRCVgQbCRtN+GlekzIfkFwaRgW5rmY665BDiqp+zkvQIG
RXFbrzhRYwPh8fZ6tIVcv752/nLLXQPVytpfTWkxHmkhaxCX+uhWwGMg4OV/fW4B5w4cnWrRA69Z
REU59fP5oLzV0br5RkpJwxgkNJGOgL/3Kk05KmdV7SeKk3tnhAu9WKVVS/P+h41GXwKKtf+xrKpK
ogxtCYYuygt+uIxRrFFUOSNhZU8Cz58nVqYZ7NH8Wvwag9gOBxDSPgbtFxWlhv5FhIWSc+syOQSv
F3ySVRRXz6seeyquLd4Wd89S8melNXu9TymIDzd2uSaWAlj9EGeCdkpgApV8g7vsiyAwtc8Zyyra
5PicBDefgBGwtqL0VvtSrReOuHWQvgDEuq2W1ydr6kivsNuVYOqIbmx8vLC+vWQDQoZI9d9OnRtZ
1RjdJKuNSz5c0rkrpRdncMiwhyil6MCsKm4NykBS0SBPSevqGTAUEZdegC4Gx/VRZNXZkrgyjuo0
vREyElQgeqfQeBsL5im1ZFhW+r4trFmYZGr0xMIDl214oq2B2mbTONDxD5bc5XOU1RDzA2Yd6jC5
al4JyC1w0xsZn8CepsobSbHQ080WwTjIRy4w+vCYf7zHy+bwPbvBmYJis5BraTpEhsYqGdT+zsIl
S5tjPd2YTF7z6vXeymJrI/Y/VBPEfJ8qHfk+iDnGDVVO1NTdHLarRr/5yAwcMRWkKRjVwEFTSQpb
8IsUaKzbaCqPW/ZwiOSw4MyNEN8yWSUMQCh4iisi5VfFVIpFyNBRcr1ooYEKngZzqHxUki+FsPuj
L5FrG5H4styzmX4X8w6CKvizEsyF9YtpxI4I/1muw9m+09Gq/nPN/lZ3ef5KI8wgpac08guBk6FT
BcDC6COWT+TkkNRWGFkbDq3qx0M5pE51dtVTKtfTLS0MxjxI2wSqnOQ00o2D4U0C36imb3se8zYy
8/qFDhYKTuuAn76/2ZqGtBjhpgz8dS/x76aWrEbpKDUyWFvZYSfWBiiLNFOuU/sjHN4eBkCVB+ya
i0sl5+l4qxRBix48RlPFhGGd5ZogYnqdftzE3yJKrtdPGyyX/ydPzxk8+6Fjt4XMAU6iZkAHQBSF
6j2VIrTfeUgOv6/+rgXdXo7mcwUYunO2iehEKYx36Rhw+VAjLT8VUKJLThMzDj0Zw0wh7b+hg9h9
EPJq2hunT6pzldseGt6Ac2H2t+T8+jQtcdnguzmG2BGDj3+Mh0an4nLTy4FlhD39538hnHS5PUku
rwaeZM+NcWS5KX9GUQqyGrKWsG5b4sm9d/k5kw6tTmIwGglYL28+6Mq8PAA73kHtjqaXrImp7ce6
KRuZR2VkrieMuvST2Rj7NzADu3yepaALSqJS4U8OR6OLZkrMKkDHusWkG5mjut8gsZokvoVc1cxP
X4nb8L4Rf4hPhAexX0qI17ld8Bmua+PkLStz4NmW8l2O+sY89zNsZR6nh/kPvBE8/PSU9VU/ZGZa
9BuOOl19qUUZD7c95hGIF9HOAS69W5uKJ7yryhNEvmkzXUu70k8ApiBZBauejwnKkUluDmiDw8mo
SEIVp0dF1mc0tynArOXTWAAMQ/4d0fgK3dZ2j57WiazSmEbga4XOEdEYo5Le3rywHQhpL12nSvTa
CPdNpQS+/o69zx5GBXEUR+GW0YTocF7n0bv/BZkdHDlWG/J7wBdRjPmEA0oWNsjLgDXZs4Gxloc1
pitH+54Mr1vszrEN33BSyInCiLRtUxtothD9sH7gTHEWww9ycJR7gEWzzLeH58UjjU+V2G2hHS9m
JCrBuU0q19bFeBnYwoQ0CPKyQkE5XduQuGuLxLUm4Dzzm2CydH2Fz18bBIN18jqL35xojFwgRRww
zoQ12LmvZsYEVQLwHfcwYwcVPaJzvlruDps03Mx42aIp6Gj1xxSCxEOSvochwnrLL4gxwcKQHw9k
9bYPxXBa1FCplCxsg43k2uf/MT6XupCyAAUeUP+h/VF7tZzBapN7vC0cauATFPYB4Yz02/mw75wp
YjvaFc6eXR+VVS8k5Qv864TqP43/GRqPhOYtxU+FGlE1F6jsJA3C+whDT9N3qOPU9vULvTqa7j/Q
4Kydnc3w5GuayNOQNWw/kIXAM9HUJCnpE6yB+TC3UCbWXIFQsnlsphI0AXzzE0vpKa0UqTnxfHBS
JcLyZlnQVWRfaWOJlRPF+tzfW2MO5Q5H51clk+vgABmbmXL0cUo+vjKDVwFHhAJnmVdfNnU+s9T9
tfxSwN8mi8RW9aQGeFfNXKaupztje0FnTxr5W6gX7Fqx4AT1UEiwRRYFaKtskEwb0XiJcC0dZDsH
lfY0r1JMOcLepnB1095wMNcJ019+cPBBK3jnB5tpvfxwTrpPYVqLC7G2UGt6Yn5iHKwf1AkhNMIN
MdlveWr+WvJZceWe6HeepPO9V4bUYCYvSCy436NYAmtMJOah631FZ5J7zuDkoZEtbFxl1k3fpIyl
rPNqgktjkqEXnt1hXYyARlQQubjizdCsP2kTSAh1JzpvRRZF5O96fqyCCIKdkyV4KTdDuOO7uAUE
lX2vbNGJSJHrt4IAEFzpLX0WHwOpOy4yafWlnVwkrv4w+6SxOKvQ0ed/J8X/E/lxd5AU1EIgudUH
jv7ab14KXkCjNnIuHQROXXYyzIiX/rKnB6raCxXGH0Iem5cq/1ozW3EvbRgn4dFKQkQKj9Go2CXS
rj/qI3f7kPOZvebkr7aSh9Mb7HalcxWbPENtsz2hc82BfoisQivw3+XCO+K2Jg0COj57pdPKWKmJ
wU4oE7iFFVbFUMv38h1PPuNzigrWgKGemG1NcK36DMth8mMrnasEDwrKoU8wSYjCarck0kElcd61
vG4UxdeCwW7rt5F8+xQZtGjHVdpDrP1wnG3ixTVj6xbwuef0jXzelrTFKLbJvRfSb3nVCXoU6/r/
8YpbKxF1PaJxXFIFwInKm+yQ95gSOSK4ggNpDqh3M3tbaG8fm60jxrgYjECJJu4LFmmcJhT9N6xU
9zEeIuxqcL0GnlntqDZqbimFtA3OcbgjkuatuH7OwQBqoPTWut6mzP+O5Tb33mh/+4Flb0j1lpYl
zTOYcmtJGcBeKTdX2hfd95Ko06gwGlZQ8RKRpg8jsMB5VHwu5IzfLFIjxERrLd1mP5c5/JRbJPHE
INIkltvlewGT5h8U9ixlvsiIxB/DWm6laDUgvO4ecgbY5fPKQI3pkWFE21KxUKuaPuL5IJu2c0Mo
DByGm0PvsnSZNdqYwHF0+07ux6nYRquDrPCwQ9n72qIyzsrN3ri0+MrIhcaHfPwkawaqLSkd957E
CgGmAhQZISZ40lqqjI3EWFH84xphJkCOqhyStGw9L+lLtPxFdnj89Xb0hO25z9e5QyC3R9WzJKJf
vlxTyPyTDIhemp3wNbupW2ilis4CniDcyOeM84mH05ruKBfssbpmPRQCFHAHDzezvzDuRbz2cPqD
KRqwyHgWb9CXuHy9rEc23EQrCIXoilsOtsk0dKl0MedPqLL4gaTZ2hNqILsITQTGR+c7xYNAJxK/
VkVVWpPMM6DfkmUZiwfqYKBdk0+tlzX1vAu7IF+QqjvNtdib1bdF1Wv/WYOLiDOCXCMCoBNDVpVA
5lKuzyF3MD0p9sLDVXauSYICkoFfnZKeHJpCYK6AEY7U/N85vgv05auF5TZ1HEBuzQnnduABMaJK
Va9yTw5FWrQOakZeUsmtwOkx7vRDfqbjFWdA9n6mevkUcB1zqHft1GNTlRYe3/cOHQ/HnbVOIyem
6fM61z2AoCP7fuJXrNiNdBMQamO6rGCbetNJiIRsez6zEySxlJPT7Sb0INewDrh5OZwCc5H9tUCI
63A8V5+R6qO90q38NWj6lqztb0CcO5a0vmSlQo1jgWaJMrhZPyR49UXs0kCQZhnCqDzCOVJJwI0u
G+O6s3ZF9VK2frIwGk+sbOQRaQMe1bdu8hE12dfIfTz6uXQzJ4qR8cHgGIThpzC8EZt+moFTH/nB
4MtNUYaYwmBu9KsVDlYYlwpUtKbYl9F8cuRcwAoR1k5N4tgRd3jcnhiQQXB9vv8I5iJnqcb8INZr
/XAKXNdAI1CI/9h6gJUtXmMtnytx+gy5bzPL8a4E306DjB6fSg/TiXjo9FrYIYn8jCjvKH4NdxSK
v7nLV3NSG8cK+tXs8PjliJnLvcRHxkAgV+eyX6a2aYmYk+cOvYleTX5vEoGIfZjPVJzhnGkxJtm2
RixeQ6OrxtzetV7OIBMJR7vuCjHQGfkvbx0L1bpRNURZaL6GqDnRSPdvdzzoCNWSsm4a4Htkb0xt
Vur99hkHI4Bm/fu0fqZjT8RuObAQ/IGxK2gRSMr/M44ZqJ7Uys0nhyaln0COf0qIODHE0cnIJWrz
yBuvekdELSyKr3eN9Zm4O1Yl6kdizlUIKfLS6VEwbx3sQWhV3CluhALVnCwzI/CQVgBvleXAMwEP
juIFJyq3WdNsRERaqTbg4NKyaqptynQ8XKI9t4xMudKhxjA6i7DT+e1TD6crKbY2kVEu6sSqwu42
vpHt9UE8WzyGwlqnPtchuZ914SwWnGBtbEvkk3rXx9MEJnSkrFf7TjB6amCZq5EJjVZgyS5Z5u6N
BL9/7EJMYT7BtUgoxG5AedgPao140j2Paif1kcybv2TBQ/fgN1RV5X+7ClUmm3cMS/cqelMk7eg/
1jtPGUupQARRKPAVTpir8nxQOgbyTtc3OytYDhyB/vGa+jl4jjWv4m/IOCAAK7RRP9VrFiYtDZud
IeBJ8y8d+fMeZe/VAbK64CM7RhajCZxZxQwDSRLfsF026yGKy8NrOniHl8WRCx1A405tjvsGF9E+
cwHn/xR9VWL8WY2HY9T4rI/PvR3hTCsPF0bNkRp+fSPyfjbj5qzU0wiSsXu3J4MBKZIjVO0nUX+p
53kN3a76o5Go5GchFIZ1N2mad8gnE0V8iR/wgqHA/G0YCjNTyeXZ9QJrdTZBbH3Qq7y2T3eiuVCs
fD0h80nbOsJLPBN+jfBT6fUwUMm89ULzU/XyQnlBpwk38SpxZIHMYzCI4PjXAVK3eg0N+SMQqtLP
gPRyfOz1vEtEaKalw3SPSBIv47hOGSv1mLIsYDgE1dJrpXvtqpQ5N24LyraOfXPYDa6pYAIDR7wa
+9G2uoltfBEYVVcjyWaXoEXsc5IwfBpYURUNgmsaDvRHoH4aMPCgUy6rm0ZXMNJeoaY7RD6hCO00
2LJ1EUn4YBiI3/HtfhsJw39OQOYWT+sJxdAwb5wZicJ7fBDBmhUas30i7JCmAQWG/a8GZTXBZ21V
+PqwrdNJLgNJRmxcmDA5gClgwca/TymkBaxpaCgytwi6OJFQXLSC9FF8FBw/zXrVNQEMlLhNyRoY
32sXeh5UaTWMWCl584OsuNxwKouZSQHCDiwqN4lQINHQ4hWqPAAJZlv64iA/HgWxCQou7kwFoMu9
yQ1E16GOIiRiwsvnFa+ze3f6TQUEi60OAjsoDxkoFgN//wP1chXTMthjYYD7iCTAMSQ7uSYxv4Vb
Y+/KHw1zsfbSZv+sTw5sko+NbV2c7XCHIHG7JT9yJL9acHos6/ivnHw/z0NXAlzcY3GlLi7TGP6a
lu/s7w0W2YkaN98xzsOpzcaL25TFbeTyq/ei8ghMdrCy1y1T8JyhsCKplYjsM+KHZ+H+gDyc//37
duApc2qD7dR/3bfruI66IAUYXlFb/uUu1Gkvv8oWmGdDI2RGieQacmmSj6RjPpyCsL075P0MFXL4
krE1/way0+YHLZX0n/8wCcJdwX1pAMIgpW7QxDlhvwjFdoAFWAaJOu6CCoFAgnr4S1Z8QnMA6TFj
WlFmTTKiR1O41J8N27om7FwTmdhmVQQBJQr0f4XNbYqaClNWeeX+VtYulJf5D8Kq4fWWVRG5DOnE
ndS+UYCT6n6LTSF4PhoeuvfaVEW/BkejqiU0tlQwvVM8Fi1BiHNRO61q36kz7P8JJFnvLpiyyTPZ
mHTOpS7D5PTFGAwPt7ylW/rBnjRgPel7FEDioXWHbNwk6R5+2nZhsqkFUXU+6Qq53aB0eS/o7+1Z
w0dk931rjZw6lQ1JBlDOZ3y/Ftnk1glhvvh5kg3y++ZtxwquGYA/wD+QtaG+ha53FIQdHUIh9+wF
6lklMVFLbv6nfBgMQll5bVdb48Pcc79JGmS8k27RpzaEiBi0Na2ZVRZdHq/SbOlYLmfnNufeoWQm
exKwBCusF4A+B3xIDSr53hdC3Uoh4N6aitrpDybmGcvjFQvBAFTIGxmRY7HxKDySUIoEL9VJVjuo
JaVVolA06euOcmunBdmg+j21wlh7do7hDGzRXcPUamEjuR6OIySbGoSuVWDGaA7NQjooAyk9czNj
Ey6Xu/24l5GVU28qtIxO5p4keGzpZZdRTEBXOUpLvxP5f1FJ+IFOAd1CgR27UOmLIfPWuCEhC/qF
7G9ARknP8Zuxn1IeDqfJy6SR1WIu9pfRs4NLD7c+tbIX13jEeNop9AHiWwYbKL6wmF3Slm9Aahkv
uCZnwva1dM8ju/UzYscjzK6h5suwKkkCAqBIiLu4D0jIaOh8QsYVbxk7IhDI5ZT4wXfmCEucjSKC
nbw4JWmZET2LBrBdAa78cQw1Oqp55wjpSJBa6mqRCEUJRNnoQIvDEo3R8qdxzUBpYPFkWkzXEyT6
kiBH6T5x7Q4u8ol/wJnXQEgpUcKZPxmYylPT6q21itTffd/DMduVCRrLX/PSmWVXlOSqKtISLZGi
KZTsFeu9FFq0Qml4ggsF9CY1X9wA8g0C/kVdxN8vFY8qKDkstm223p5g8oybJjXre1pYhZrdDpxX
cDBZQNPbU881Kg3drORdvj0VkqXSu7GSjEJYVPqaP2KELK/LRFvlEqWf54/KwYZ8hBKELSdFf7x6
qZlIebOIMvJw7NhUbimpBGeRjSqSAxxmf9eifIDXbCzRa/kaafaIeykDsu2iDC5GtQuJ4Vdr4cyl
fypzE3kL0XLIPszRbgYZWDGwEv2nmo8J7X9FS5rDo7Bz0eJZNE6lgJ5In8xC0pkdN89DppVpAYhE
BggTfpTtNKTOa1GNVuJToQodxv5rU7vDzz8dz1OSnM/YW7UGazGXurQYh42GUljRaqNytwohJbw/
DySQ5qpTxEVqaRDPwNJC0X8FC0rRN1p4edsMRnPeKVDldBmN0h0hSxEqvi1Yxo9vVULn4LBnNEAk
gYZ4NA70RTvtf804bxhP6YLSEEOlOxmdSlQkFOKnamozl1Y4x4WMMuK+UTjEPaDieRoXyw7xKgWb
XKkt7vvGZpb7eGvmchP0g8algtf5cdxCLLiYsH6V1dvBtvRwkWy77tgrLuCmUs7d2PcU/cY2DRgU
0XK+wAshz2LJYmMBnsx+bwB0bWs9n/r59l2d9lnK6kwSqtWuoFJXBV5ujxBbe+8j+qDY6HYY81QM
q92/jqqlFBMP6wynGY4pXp+ArQvwA/sKSUSrOSXDbIbgbjCZeGV6sHKWfq4qL6gHLOKPsD+J/IzR
NGRy3Itu7pZ2mjFdaOs2dqdsFeE+KbzzR1RYSKnURxY/e/K7oPLEGIfoNaObwQRGjk6ngCH5NU8q
trQ8wU0qhLzGZoBnDd4BvaHbwSpGh10wrJqNMTAAKYQKrTlM+aLrntUaBBDPuOifPl7QQ55o6S4Y
2qRSiDlR5Mz+2ScqNX+M2Bq3AuTreOqydbSSvdwD1wypC+SwMpbVpfBeaeVoQESoEZM6SzL84v/g
ycpHhpaP4b88XpgfG6AQ9+oyVjZ3aUTD4m/k2cm8SB2nkhAx+gF7szcBA+wgSMwKrktAyCzH6QNs
TQ6DBiisB5Gm6S4CFvNcb8jUkTa217/9uHMOJom0/1fwVBWMzk53B5ZTUl4ReciQ0dWdI1AOY9gw
6YYoCpxnurmyiR4K82cp63NDKEVbwW6HrYsDWn3uJX/DGYdodNSHh+GBgPhRvmuWNq1Xn8U/ohbz
KHwQLntesyCEbxrHrkeNjP02zEirwdzFME6tEAJ6mHBH385cILhgYdYXRMjLUY6ZabUsc8uOwVj6
mkD3WdVrIuawmtVmZ/gOhh9weK8eAixxakUuEnysugp9p+Z53a6cMB/kYMz0pe2lwsOneT/TMvKQ
DzdT1Uj9ewbwXV33ySRx8UTA9heuN8GNSEfQ2849j55Mv+CEvyXPtt1lMDoV9/1pd3V8WIilr7Yn
Ft3Q0p/uMYWPmUB4GOcbEFzNGvr+PvQkaj3uIyO85JfFv2kPqGKG+b66eOg1XvutK2gLDYTwM8IF
g6kRxQJ4tnkyGlwq5nYLvhaE89bMoEnLf65QNClrshwilX9FLP98HWyMFWYVT1BsN+PAYxsa3HtU
fZ5RRcUZGGpNd9/SchrFsHVVRcLK+5jrx1wCEqE/rz4ZS0I/FNyP/EgusTRGjaqXO5v7zfdKhzC/
W0sZuD82/OKjNZKQGqKW1oxAuT2f4L/T9AAbgqxJZ+bMi0IPY87rU5pV0h/ZMPOvw7GZJEtKMXs0
/7+aAcPpeKsmsI63DNs59aywAWklPKORbJqJST76d9BALbt3giO8jEbR3H2zB/80DOe7DG38H3Aq
2He5JKjkMLYgXt22r+PGMiEySUYFVgWx1KWM3wFyOB0wlOPoExNgm80bvi0Y2128emai3u4clN7D
gVj4/TFG1AKdoQo4jzra6QqrsQ+xzllxiIUk3Po6SbGPl9BZdtdUXa4tYGTtwLIFRkOavddynlCR
wTzurNfPaIQ3cjgY3HeHLRB728/o0EsKwNO3mCUZd1+ljkaMB3PfdNH4KCNXzWGpLcjF4ml+qn8v
/fUCeKCzSjhtRJORMzdVhjj4L9EuBxSq1UQzwg3Q3SMkGn7lkXT3IYxSOs+9Ap1gtDHojuGArtqo
VQQemACBVVIPuctmRluSd/rt8LhLGNxKxjgj6bFun/msaBNc7dK4lumA4JFRQpOLfwqCNmSGlC1I
qmh4cW7lv1ndcxNIKc6RpN6RQlh1z0CQG4RaHvDuNncO025heB9UpR1uAotd8kWWLOSjQ4pwsp+a
eaCnhYNTzg51tyyjP0x7pX85gD8Z+TP1ZmrbmsUjK5Rx9u7mxpVgWZTFFeuk+xtsUruVdRWGLvVP
8VySwl60hcuWionaJIP0MiDxt/gEpV9Tnjel3vDTKdfY3qoRVnUa8HIfZ0rM38zFuNc8/1ONx91j
htgwBbvlPJ2f4AbdcEBmvQ2aWP+Tst09/sA2hmWCEni1Wd1yZvGFqySdkFoM2OosLCZm8Hh35VP2
6e87fxg3+qcHAHDmPvmqQhFBje4mikq+SyqyV27LJNahTKCRygvIF7HXSpyyZm1hWWO4QXBy5+w/
8hUi1taOiG+3MH8mT6mD1hRgTbUUwlJndhSGhrPr7Diu0p1IIEf17lLtpxqGE9TrUal9cMwYDiuC
HfboL63Vt0A8KkDZH5IOgUEcikUNolfTzsh3k4L73xn+7XFjCxhNivndRMnIwd/BVdWoEID8swEY
5zeIR8igtetQ4evjULIbsmeLB1D3bI23Sl3nfFizBuF3uaBm2Bt1aTfH6Jf0gDyaij2yGBILoDKk
5h45fzMyBrknPwIGyMx5syZ+0/QCt2YjIDdfvGMufzRvggUzWeOa7X7u5vDj71LbW9ZTHnUNhiwD
78eUsZ14Nke8bQfZVWcMtFLyE7ggqivGz8D+GQdK45SyJoHwl6db76kXWdwt7tOea/FeCTGDXmfU
3Ee0uZO1XLh8VgEFKquTgpWAQtgpDMYK5ziXbW667aMhb4IboeVuOd7ccCExxs9wkxKjNQT05Eks
v2CC9EiMdpybijIMexKw9gUsNlePIw4D6Vzw0mFdQx0lkAQZKkiuezCm+UaJ8vuSofNI8y/hLng6
xZwBdMEbup4HyjM9OS+o/dhWpmYLfe953JrejL2+BNuer/nFhRzjsIs9byB0iLnIYKhETKR9xDRX
ALHapud8QTVTczr1IYy0c8WEj1atB0ToD0DNxQ1YQJ3gOrCiUNOZYlOSnKh0mEFmfk8CSEgoEvfO
nGeNzZfZMfCDFmS2zE2vp2S4UCUiQmON5amJdNmvvgeVVmiIVIOcdZUGvcEhaIMTON6raBSPXr+C
5HyFvrtV2unH2zNuOZIcf0QOBNU9DPOw/GgSyWKMlFMrXwvWDrfClAkUp5YKX8sBV6ej2sH95fYl
tnYU2VfgFlMaz2uJ/sDftL919NPqQVaIR6RVCcBu2tQczbkGLEjMg57YfNkhEDaMcaK1KsmG5hOp
1kG8EjbVv0t4qdosMZNFJenF2XOfWogU3ZqQkFJCZrwHLmmwu4oiykwLxzw70DbtdkhnW6BVo13l
Dyuls0SdY+1O1vFR9DS45KeWBCVmRXAN+kmcT+890ali+/Zc8FBMd1Zt1GLTRQsZHsS9A7VjrqpC
tNeDq+y/ohS2dr0hHXccrPa9ADkPrKgjr2HHVqwCfCyI34Plwxt94+1GTQpTXVQgM+ETOa541Qy/
MSeHQpyjzPA1Keng8suxb+yMU3trJ7a/GliVtkB7Dk8P8xglvrnFczdKozU5Zu4ae+DTq45QaHNO
zCsNgXPrjxA0YCixfeUDJbpSzd4XYzhrnk8LAQrLv6Ndk1w0YG+KpHK234krhX75pfzoeL11HxoT
U8bzQW5/4SrXII9CiJPU9aceuXVqg1atmLw1n1oML729RYPfiOEK9mhRR2bFrlMdsBRvrOatNtBI
vMb6CHj5zjPehyV0K5GZx3kEB291AwfF1UU8R1NWQJAMpRjqxkfahAVgZ+kVI57WrPe4PMYx0ZTa
+brboxRA9QSPonv4Pnvk475eI+wrxjdqh84r1KfCIr5DE/p25LisvB4LXZhja9xv5Nppc+bGvLA9
sENSFpQpWPPjtds+wvVVBDNjRxmOl2C0cQDkZcS9NGZkOyZagGE1InqUdd6+ZJMMSthIwCCDel3u
73WOqASJoadW7v5XLzIVrnW0u+tfdMOrP5ROrt+4a+WWyUMd+Km+gysKU1D53VM64Cb/wGhhDBcQ
GMkcbhhtkWwj4ae3jiKXTgjOoFnefUG5J/AdCpvb+f4bHuSY8vQwRbPnPTtEbpctwKvBbuqcgKem
KLEstepfU8uhIX6hUYNRxAPPsXpJj16EyQR25gK33/nPXScO/btcB2mSB+MDdXD/6qAQTboKh3B1
WVZjl9euL5F9Bb+Gnwnu+x/BGxGnBRnPIzKeYO5PrLjh9HvsswMwz6tJ10ehxHMi3SeSODf3bWDT
ZoG1afx0wqF5rY7P4y6CTy26yr9U5YcmxbngurR4D8QkY/JX0xAG/uA/GhUS3953/uLR7ztMl6HG
RHJO1VPdOM9FDKnGwu5EssP/eWf3y2QBKmaJNB9bf+2wulH2YTFV5OiiJq1PiIjs4zbzgRZirjN7
3kHVBRmLdqxpzsjxBkV6iaY1qy7aHjLYnwChYQAvku9JGZPO8E1di+tqGcma6zmMPnjm+SPDVQ+1
ZusbIQxWHUynTela7fMiO79fDhoHi9ivl8yK/UfJdH6Oo/V/y5ON6u4QGC417KoxU/oxxwpgJA9P
1A5dFxJIY8Y8VMxj4wxxINxVe9arvm2bLZML0T5iJ0HSB5If9ecCi8mwUhURL75L5alF6UwXPFwa
iihJ+TEGAD6G3F2jfElvlAYbyD/C0hylU2RjRoe9D+VLvtL1Jo9IM627grzUYXBkEkxa6mf5gAPv
Kcq8Uw3ZvTd1pW43hkvxVwDTc5+oZ7XFAlXtCgdsnDECT8zH0wjVsfMRGHygGNUaW4EoBNKpfTIT
uRuC8b4JRukBbAOySfSnm5NKYZrdfwwMOMV6xMSU+XEv7mca9nT+S2NisYUJ/SjOWypjcNXgJUMe
g5DxW9WtA4BQb+6XkuV1UsMSR3du102kq9wxQBU9HdweZMrKSJ+xnLGupkEqPXPaGTUlsm+81Au0
Ejn4UVtQx3r82qyXsB3n/26axx1uVToMPX9EMyiWnfkX3K+OPBi7cjDU5C7uafUuKbAiVIys0/oa
FtabDQPleXxnmXakmbWW8bLn7yDv4/VE1dxl2LpAvMVh46AVwRe9SpDzwxVAkLqLSTSvhdOKGNvW
X1rcFOaNDTJtmRAZMLCP10zT68PE+g6ZSzr0s/aSftHDL8uKLj6LJheTecz4GXmi6A53TGnd1uK4
mjE8Xv8vjsOrRZ/Y/BX9KyR/KevLBHvk0FhYtu5Cd+JK4I16ls3WvO+pe7cIxApCPQGsmepr92lo
JHtHE5gPcdHsenyaem+Z/LLHRKWhAwd7SFUqnsdqMIAwYOaV/lEnm4G+dSKRFVacDNp9NJ6LTYA+
ziZpdz8doA4SMpxGets6mN6Ej3Rf+nrqAIxoNT2gznrowPdkZ6CqzOoPUZEDF970Tr1ohV0PsERE
QcQJzwt6cvdVx774lgMFqga7SLSKIzoAkOXI0YFRnlgHhFOAn76k8gEXSRepariZhcDUqErfLMFD
L42c0fgJP7jiqYZVTq86MzKtIWS2QW62WGvISYT6JP7meDo9CTxGDGrskY4LbPsg6i8Uxv1CG0Gn
EtXzXlr1BiSvXNq5O31D2LWLNPlNt/myVOkNRi9MsQz3M7lTmaONMM0QZUWBMyuj7Y4Tuc/pNPlq
T2P4wU+d/4TtYjlHyOjVWvct4Q/05tV/j9PMar7nrw5iQn0Ra+l1Ht4YmDHW0ls6cyY2Rxz7++tm
dVwYrsl1EKxRZrPsQ823EVPqfbUJBcs/GWyFmMMi3j8ExX3At6mfZzf8jv88IXgF91a6fKjpNU42
Cqg6LMUUf+MI+mWZek8waL/KARPUVgJGOapCdrx756Z97I9wFgEbBhPMjufuwyC6929GKX8LfXF1
cZ9CEOXZ2lVyvpytqd6FD4kzSlK6vIKt/V1JASzIFNkV0Y/cx2WUmgms8rGzO79wDLQ5NQqXZXwn
SiGv7VYcd+71fSqrlc1FXUgXAWaBh01E1z6VwQRv3ZtHRPdSul0x83AXxanmUIC7u7fKrp3uaiWI
3B6A2KbaTIxG1BF4Sfbyk6Hz7S93VvhQ+6AvW/Wi4X6k9yqbKXKofdCXQ0pLWvouXylg/t/f6G9H
6Oq54Ih26ejhdD5FlRTAVJWg27jbInqTP27EkTVaXAChjlFy5C3vNklSDXz4FcK1TrekI/YIDYYU
QXMnUFLeGBRzvVDAz1q5r1ZqkrHO1eruHcHZ3tCCSEBInJO4OMPjbK3YnMzMN9gRhaGjFZ8YXXzT
vXB3WBpmSmXYPcC2dTNW+i3HoGDDKMk5y/hwxpXbqrJmRrYKUD0rPSYiRIHwMNNa9tnEHp1iGV5T
4xk+rDkc0xMOmSOjUvEB2XeXQSVtjpsnjrX7nPoygqkNGaLeODYJHgTyAKOfyo62lKwDRwnWpFvy
eS+APbHY7vCbqH7p5jEe/YnQvcbO+uKG1GUUCm80yfvFLveCG6AnzOLwhsqeEXwdaG+NzRlHms8B
VHUe8xWx5CtgtAbTsQRa7vPydv7Bj5rCWwScLf7nikkpZjHQVrXZwDNI92gNRPMJMcV0u4pRvXCa
AAsUu2xN665Aw0OmdExSTxfE34NJKBaT2xUr3kRtTIB01tIi1pnuKw+X/qBzvfgx+XGcWeyM3JoG
+/z/VDigTHcl4mXnrHmvTWbDtTtNjzWTRlkyB1pFuX5iSdTNBjN84JCOCvZbX8eebiv8e5Ot1oDV
vvQu6ozNEPaj7RmnoNOXK7hDpjRkvJQDqJlzUGO0SpH0e/lQ9LtNt59XZBgpNwDqfquZVkL2j/Rg
Jv1zykk0Z9k337MIRLA3QBl4KXtqK+QnPvBxqsrMB4h7TAOFHltysMuA866BMIYOtXCCJr63wC7E
nRmptqDOJfZYvkSd8J6MYfrHTyAwvcOasWQs3JRs+IUvPIufFkkVOV+etaS71lZvFBLvxb915LyF
5MrqYtlXfBbLflvuwVrrW3B7HgcEM3Gs3GhyD4rB/yZNsdPt1LkG3QJlHG9eWMNHoUtkzOo7JE5R
LvWWMdXIPq4U/5tXB29Q40lxIGkKm+xQkjqBBU/PkGLnH2ptKrdXrDKKBx1GlafIESBaRJPeFEio
e3SOFqR6MHUZtQhASNEMLonSW1eksLatTVYczsuMjNZQnj3CCLzKi7amOg8JHqboUzZrcBvgqXeJ
m7QScDvgFtgafWfIfv0NJ1NHs/LO0TBRYFvSdhV7FcTdPqrA7WDnshBQiQoFNFtA4eOrooGn9Apw
iaZKTEkdxFxEr8few6DRHr0unbZsO0y8pe+dpi2UAlGyri8QNsJnoVPfgjUgjqB85h7pBlu81QKE
90peCOwjZcqzU7z5o8HfSOoGKh1tjUtHIuSYenu4uhTSj2Z9lT1JB5Jvv7V4aAU4aGU2tturbBFv
pnXtkm7ZCMR44WCLbChHyQjwM0W9yydb3Zd1oclgdvYQRJiZxrsKsiorqpmUTDc7pqejToYkqiy+
0P9kUttbSyI6jlCIeYPUE84UH/5bTcYySVg01pK9l3zh8xUCvZQR4eLs8Qts1CItVMQFKdfliFwk
VZW4lBneycARq7OfG1jj7/UOY0KNGwNdIr7rwnNMy1/nulogSu6LVnpu88UphEgBKGAN8BVKrAVz
NrjfzXpomGVPVrYFghEosWNKS1jCB1iGjhh4NF4MmYc7h4HwDVto0LgyJz4Tz2KaWy3pWFMYEerK
zRIlrkLOCcOWpZUSLPcYmJH4FbWXfANsfXQVLPBXFPMqi9QNvjF+z5kNtQUfFhp7Vux+5FrRnfh6
Nb5dsMw7HolRs1Ge5oUlp+bP1zEUA/5goiYX0lVoDBjiyx+m/2xEZkjc72yxsHcJicSJvKW8C97j
Yzt8YkFMPO8A++W/DHf8tdIW5fSLVy7Hbq4UTxluRYdzpF6y/GnCj/LQ40O2Kr/gjwdJ25dPr3sb
uqXBCwsPcm/bXxfhshJAwwyXjibucWhO6sKQR5RoycdFp7YYLuADoIUkSaD1zLuVUirI6Q9zYcrz
grev+4NktINLdfazdpnIU8yt2vvV1pBVp3uTq5VVhxDG0Fcjg5tPi/KpdDXBSk2OX+14E1tkbtcT
Ca2d+HslCu37y/WQ+OcFJ77668gztgV0LljTt7WRaPhmb7TsxS/0lZWqYc31l5j0DvvfQwqhBCxR
gN4/07nQVMJpL0rZh9h14p6MsRF7HIVl7gbCjJmTyqCPT6wbTR3G5X76qD+ZOkgaJUqQExo+5bgD
9+8KlWr9iNsm1ST0U7AvcFag8b4bo+zUrAJCTMgdxFPS4DmcFJP9CAid874UypFHGaBReAZsNnzu
5oGpjGni7GkI34F+JT26GboV7Zh7qkrB9gBTo+MZcplSbcPpOk2ybcihLPYCy2/4l++V1eQurs9m
nLFZjlkVc7l4ILfySehgjuRhwundVEveCWzvQnYtBtcNdTz9etTYXT17iTz1L9/vZ/tj5UNmDWhq
s6Nu1oNT2zEFHsk/L3DqZ6tN8oqLpJqdj8/fdUbxUWqwVR6dXn4A5kEvNksgcJ7c0u3kTtsSpqp8
ypFMVAaETszHOGIGdr/tUS0GCbvNEtH/QQcbI524uzGiQ51eYs7QSxCK+yH24lyYBANiXoi2mbBx
DBjltL+NsYdTcGtYv3rFpnc4fN73K6GjvscdrTFuxQ3/e1TqR68DlPVnFMeyqOo3y6lMBb2Ne6lS
wQgWwoD1hbOBhhE9IjD90LKzIEcunqaNo8MU9jq9c8m98QVB+2cVx+JXvBYxLoyLZp4/prX006af
/K5AT25aSczjrBs1ygGM1+mtYMwtDHY5100ZRP+2zy46znp+glSzopHBuQVdIhNBQanV0px5GWNI
DlsXv2m7zXolDhc2wiACqg3JoRu1VrpK2CW54lEbpx+K1asRDJXquD9w7HJrOiMNb3rWuexu4LF9
DzRr1MTnoZiAoc/7HefukD/E2WqGASUDFbNSQGb99+ck1nfnCEB3vaUNPMuwncxa31HNxfLF6jHX
m6W496iWEMQOV/iv5v0HMzdQ6oId+M7GRU8vHOR//5lyOfkDliEezFHjQ9+E3FFYSP57kPKigKvO
MCh1s0DKIKvueMYpcWBjeT7lcmZnWy8rIIAwj2YEvKQf/B3+YmCCNdJbTjGeRQwoP13QH/rfABwc
57Xs2rXjizvVic3Xv4ySCC21Fp8sTBDIcc9r1tEHgBrt2xPZUGBYaMuBi4rYkhJXm6hUX31SSu8C
dqEo6p7UqRN9Paj1k1yeSpxkDTfKSzYSeI3ln0Mv2ilVzrkXSFHpkDwRy7nySHA9Rlw6XoLm+Auh
jwVPgnPFEc6uxxde1m0I5JDrFCZVSa+bc23u6fTN6AY/MiWGmXaY2Lly7qTjxWJrV8ZvgH0WQUVn
MYQyKLtYmAWzcuMSHywjCzrAFsTAZEzs4D1dD0P2ABjUhIq0l3KVTKA5/wciBPiIdz4NNpH6FWnu
zzSZ6q/FIIcH3Mg8rFKCJZqZ4p79VhvgBCqZ+lA/FuIHPqIy1UQ4MXEUKgWQJXr7m6ZXIke0CZuH
a4ZxKHlv4angWueA/6QWJbIqBaAzZkD6LG+6XSjU+SZ883kVdg+mUazuWMKbL8a5lhNj1KkxsAMb
qookQBjY9Yh2LBxrVuRxDmsQBmRTZpzpSGcfuBSJ48+qVxl90u4j2FR6YbpkeNNO8U5BmiCFerGC
a9UGqvBioon2wNEDbr+Eze85A/mEw1sthRUTgShOz1HY7IjAOVMgRD+A0E7aBa1Cb97bC0KTjJ9e
ybj8edwnZm7JjSSVzMeC8iYjpejjs9HigwSUkb0I430Q5WlkdY49NtvxKaTgGUR/T0lj7pmyVpuV
1JKIZR2Nnamxad3KIHhxIH8R6ZXvnDSET86SFHVc0xyeMCpiAVHqotY3uw+yU6TL5fxb2aog74i2
2uxfJumjGTaHk4fQW14Pv+XNs3H0cMXAlOEZ3kmcGUyhg/t1/IeVHCubRjrUgzv9tZTdf7It3dLz
ZLhplRnJSbsm7Sqn5uPvha95p/46H/SipN7xSAR1Rr3BojldnB3J6vYGQTCblACKNDlkrVtfB+Qx
kcP33V3w9OsD+9AqzCZuWsLEmOp4UazOaNOnsUYm/HT8bJnZstpvzmZeE8uJwkGuE/9feFdhn2cU
IAi8XQaHR5d1HOyW9uF+U1i9FlVQ0B1eMvSf0mI7Dh7nm3oXNTrrP3FEXq/7DzTnZ9c3Jx8pHYSa
gxQnq7afO/sf/sjo1YvNCghebnFyivtSVphRj0PCiGiLm3kuzxqydvdkrO0hR2q/zqr/vLruo6x7
1PypYsCXb0mzexWvC3fEIgX+GhrWv4HpGxGwJbrqZiOwJbvy5MY6sknfrc5ZdAqtoZk4LwmRlByO
lFcy4IPBHoXELTkYcvHWsOKa9WKEM2xnJNuK+s4CA0pBKs+8LX4GJw+cst/tey1Yp9PwSPbUrboM
fvu+rv+826Jl6Uxf5DFg2eta/ZoiXxVOqM/iTZvaagg7AQtucyDAnVdbHbnjcZhCh86Ytl7RjG3M
O7p9txkj77ExnLWkspUkTZHg53fbKPUsdxhluGWswQpfzo6MecuqCj0Sn/twqgpg6xrPgczGJuzT
L2aAQi2t9GfLFtL1B6f/Twk2UqnhRF514P1OYwbJiFTNfeEGkePocqgy3dd7t1CHwc1JZBksYxsQ
j3OUJvkzcmGYOKJUK9pEtXyxHHvhoQOnEcQA2GZKWRgqPBVGkbhPJ5RzXt5XCMvunGy5MKSqnjqS
k9aUNNSwIDVRkbeFXCMcfOulfGS1vW9lHBSXYYyAXkX0f1EK+AnI4Gp2q0uH6ov5EPXbPsI05O6D
iaVOzrIVQzQXVAeXv3iw0zmSJi8voP9ZLaR0NKs7TrEkjwte3E+j8NUHbNjKDNZQT3mqQsR9zbeH
mWvWCcRGUaLSxvx6IIB73vEq+8vn/PC8hjSSHVZ3yPZ5/DsBqKpIVlzUR3NlS67C6nM1SpmMu5Dp
prGIaS/LI+gOLkBnwj/8siyflq/MeJZ9R7uz+YmE7NnzdXhPySFAZb6j6pcBakrMDzbFmEbri+N+
RLFIkkNjRTbykblyleLFgISKrguDQVsDYTrD+Vjk/2QG0Jt6682FeG1FrH7xevla1K3VI2k/2IKy
MfDAhMXvlowTx7PK0PinRsu5AT9KTMGO/Bk4EIssVxHCtoGSiTnbcpPKQezPd8W+oG0BsKQ6Qwct
+QpIv2I6h8l9/7Z9iLg3c1Ax5M/KUkMTOYg3gMBdoC4RBDkHLHE5oX1N0/uQVljEVVSdx5TLwMUm
8GBjhVVKdBya2YOyPwO+lTylWsb4lZEK809wITFSoW0YLl+9EPFMCpp0moZBaj5s8d2+CaQQlh9O
bmk1WI3vLG3naatCzy4JKLXV13IVA3EDVYnc5KA5SmXdf6xZUV3uhneAGp2hp9VxjHWNlSy3tRQz
ShkZH27vDSg3pZttV19PhGkhduxegJrRr4jrFfQaZ1m4D8435ChLmTrOV+6neGtNEYOypFcxlR7e
PNaJ1o1qc8dRFDrmR3Deebf1Xsbokv+XFj2TL/VFu3GMslhuAAG45konYsP1nlMU21jNjeDQY+fe
nhx8a/Nfz798z78NRVEnIMYrLz7+6qSCV1xc/DFR+syy+blTC2JifK+KS/BkaIMlu6UOr0dZ44nE
0fB9V5yhPXscf7MNo4C2YiZW3N+IbQwLcCgATJ5zkku3EQAioEbibzj6LzwUe/zsG46jJTlv5sup
zZq4iLcpDr//OV2MEP9vgPwqPywLC+yM1eK1shxzaUjVw1AJpm1p1t2AJDwKYMlFVgmKqKQ9st0k
1YpIu5lH16ZyYBjyxD8AVs1/rWKaRE/yMRFzofGFl706AhKXlbKYUdypOEm7cRkj+0lSZL5kdagp
RevHTVph2C6F0XqkrdKlmsHYJdyoyJH9wXrDLqoksEsoCOIrKC0ruia13T+J9NWYmsrnvB6ZAOsz
E4NbVgTL6WtuqqGcF9rpxKyyVgkyh0onS6j8sy7d/eWLXafjnEoYQ1FG/4QpyxR3CbMbgqx74nno
3UM/tVaypQwLVKB1MxUlMHXQVdWcgvMvUhJOlLfL3kttRHWeftmmdkLC6jcnKLnV47pq34pPeWiN
8n5W8nkhkq96FgjFQp5Fy5xRIIKP0tGC9WKM8GFOQYgGbUcgCJ6BQjbXUypP09/OKQf+IL4ZzMrz
mJ0IUzbdXhi38Jmp/lhkWQ3l51xYgywHSome31LxRAmXU3DSz3tZ8F6dkS1Av8eOj8E87dWHxGhM
6yUop+6JeQCzg7M2qT+vMYQ8u6wZ0TPs5ubUEqcvGP1Y2KxO/xiLJ5Cj+HUuaDOaAMC/YlSDBwvq
Xs93TgXMHnJ/KD0J48RlxVV0IUFAMr/lAAlVqgQFqo1KXO3Q/cIVZ+hC11jmQciAvk3mi4l0hx9P
BCc2mtP4tYVlKZyMyBPHqsDC/mVXgEBTXCA6Am0g5pt4FoBjM2vxm0NjcpwRmqk9my+A2YC2HOjG
lMb8sUBGm9pGeZaml/yB2jYRZhaR5z5vJXB0EkZyD8YJFxbxV2amnGgEXf4vaciQ8nkplkJ0Cwsn
bkGUMGZiJ68YjpXp24vz3Qk0xXJHceyIypXpxuBVBLzkQTSkweuxoAQ5N8hsDNLQjCkFQ9UBQFZA
6T6JzJHbLqD5e0l+CI4p+oPeaXzp/VMB6b6yWGQqOmcmVDe2hLH2BB8O4x5AXssxhtfWi1TD0AMb
9n+XxnCbRW2u8/qQ7E6GFJhhG/aCFFG19hGpAnGifYX/i7YVIVGaV5wlh2vcUV90FahViR4Jv2DK
Tt3O/BG2PKKIzpqD/x8pSixyKGDpzoNt7tO8S6OaLhVHE0L2yNngvZx3A4JWdqwQpt9AnN9P/AxR
UQDyauYr+h/1IN+m0B4Pr5bO49Flo5slCdOQmS9+q8uqZlD2Db+0JxMt+ytYlmyUcS4El+9aBQji
jZcbxzT5Dk/jbIRcg5X7PUFlkWi93i4DfT9iH/CzP3d69+4Hpyujfws15JW6PNtvgjXNtBrRxYgT
tsckOdu5YWFds4G0YtL9D4VkiKSqXEbLM1ZtlGvlhgS8AWx+tSnVOCau3CD33zdxhQ9oxzEu3HQm
LGGAU6l2SUWOMfiGmbRKRUhtK17xVvm3nItB743x2JPYot74ubQvKA7YNRedAhCt1j/sViI8PH/x
CBdnqLyRDrmDLFryfVNyW2yiSOL2uuyHwgjYXqT+4kCI3rRQmkcGcUkCCUhrtyp5ih05L7+cTYa0
l821PHenQmxDKDS68IIJfum1snALRIdsPmjfQaOPInkyIqFhW3gS7hJ/3yt5nR70gEKMcIbQQeQg
pe5AHJJXlvQ1/y3TnLhLv2LpXCoA+gQTkXpB5z300UZQFZQPv7pPjEfoHj903f6DWviO0hF51qlX
B8drd0QtT2Yr5kkm4JGhzWfOvm2PYJ0J7dxYZ9DSpCqhM4UdGJWWELFDiShDCRG690OwTmY9gWms
/fyciwvG1wHfDAE8vxN2HyRvY9CEOQirffM4rscdeEs/psJHy0FpjWHbw0jrcqXIu0F528Ltt6nq
KGhwpy8A11OrtLu2ZKU6P1ya3ZvvUUYs6pevi/loqruOAcqS/uPkHi4ADNQtPq3UXvhQBXe7El4z
GSZIeZ8O4yGWjYYARNKMcY+FGTspNaM1mCJTpTSmJF2AdmuIXlgL1tQ4VNZMa6dWblUkjUk3Yp77
HF3qrKhCLBC3v/DYgKh+RtCoAV5vwxZzAGOfi+L1YUof/Fe+JoOC4E0rzl9+D4n1J720TUuOTLIs
tlTpmb0stKpI6SMnMj2kiQIa0PLxPWsrw94kYViBJfVhR5hoF+y1XJ9rbylShR8rd1+iBjbDH7so
dluevzuqHh0GQVyIVA4Q4eGXegGnhCK2IZ5ywncTnHji+wE60oz3BE1CNubteZ8zH3/IuLcnL028
BWAtD8AJay8aKrR9EqYOOE4jXUIzeOpuzlq0FTC1MSpaty0qXsgtksudHitzWo6bkprr5K7UUo4c
J0p/lzj3+r5jcnpq6mrsIycudF6iXoBPFPpqEgHA4YWGxRqF/0VABnFCnAZRflvntVJ/ET8yC93K
yAbW2OXS5gpjEtBKSCEOQD/n7C8TfCaheYOY4goHu3lDXvh3LJJo/cEe+BWxEMBXmbq/nAMXOtFb
+V5K33u6K956JTGu4aBz1SA/0gx7aTuWG8REt01Ba9aqOMa4DUetTDhbMTbE1eivCZOAclwL2K+s
KrI2DbrKRSXqmMq346yFLtgu6r1KmUZcxwhytZHjT1I1wRwoyGkM8Z+XdjR7GUhmCPN+YeIms4RQ
2y94yVx73xgDtyqFDEYLnu5UK9E7zNEPEhnGUcNToM9Zsazs7zDmu7OL6EVRZ7PI4dhgjTJacvYF
AhKIYomzl9/pV3ZETkGeXRgye5CuSb2gX9TuVOq7TnxQx8gzx2b+BT4JFyo2sY3DsUdzgfOqy3fd
Kb6u6IksncpD9AisqSU4R1VbSa8EmOZTGbTJuhptiJpf0ZM7/RoRFQ85ySjDEVSvBxdHUQq8undu
bBQEd/vBvhAspkP+okyyrUrIwrFU1hppbYm3E08mDhfUgD6X9lccTOqSqwnXJVe3JHUH2NMHd4rP
bYc9kmTGVAvxlSEusoF1F8SxgtDIrzoxi2A9UklU6HRSljwaC6+hxAOSCK/XF4APsQK6icS7Ux0A
LNoY4Tz4c39qkU96QyKolp+4jySwBNhx1ECpCfkLVZDuewAM72x+SCD1oz97G9+0SQTzR4pKuvSS
y3e2cndjIznaXr8TmWXn2Xl+wbjLMkiMMsvFRWeYiClRHpFvkInN6Vb/hyFOYAm8IB2b9cA+lHMA
abJSitgq0TtSabnLFqCFbk+A+l9BgGVrmF20GAxabJTRMHuGSyf1W8LjO7CimUeFWnRUcs6+0IcN
0MRYXnldFhLYc0NVnjKixZTp+5tUVTFZZPSSbA4TZdnN3yusYxLh1PO1/HgHxazH6eoVt07RqaC0
ebxW93zwXCVLjJNbtTxXle7ViinP8Vur3QiQhhAZHmNOdwT3QuG/l8HmwdKPfDf9jMAgUyH9CJxh
cBODjmZnp7OraA8E0JHufi5ima3QuhQmZUZDIOj3aWNHlcgt/Rd38x1IWKLwMkJmNIAlGLcb81P/
0iGmWeLNlwZepky20p3S89Epenfbebsq5jUvGxqksUeriJ6c0MqhhPyEcjLjAFMDCPQPZ1kp6Ty1
d0FiFq4g0RVUIIE7LQxBDYepVI/OuAYPOzUcS7d1IW2uq24iIaRFQBZar0gIY70G5OiT+g+qKkdJ
No4KHshRW7ePwv6IckjzrDpKdyOtQnTQCOauQXrmMxxVIXtzuZTmhqFYORllCOlDnY8z/6nHV74i
gTeZZ38TSAxz68huSOYOwCSevyEfGdD+OTsDdBgHvY7J1N68mTk8LJgCy7uQluQm/Jwhuh8SCwWR
nBZ3Y8GsXy9+d8Hm9s2QPn4qwW0EN1A3TG6q2lSoFjuvcN2H0kZToewve/TFt24A6UC05//z4ofs
YEss6IvkoLcIsxvmi9c9SSivoghes6vobfx2hbgMTLhjjO4JGttL/vesmSEGq6rONl96GUZxlFoO
MQrz4BT8Kg9LB9meNX3lEOk/HyIlZPMRF7eTM2GGC5xgClWSvOcSCpoBX0vchOlSfJuZE75v6veR
FcpPWXtAmZ2rWhIHsEiIMOHwpVp5ei+vbfTADeSmmiz4+ua8PRy01I8zgPO0FJl7SKPTmFKh6sDW
yapBWPWT8sV9Fm9ihUj/Pxv5EHspxt+n8J7n3MFLxXNqu9CYquWZPY6SYVaEAq832JpqBBkpsFuT
7FNqw68uh63va4u1eC01KXFMCsmm8g/3DiS3yZu/c9wXYkcTAYCUI1wNQO3FtMXl66tOsITJ9sy7
vtHztCNAJlubcU/2qlx8/tmQ1P+7C74qouKwU6lg1KTL6g4dbYvuSwe27L8//fSZBVYBh3XukLme
RwfKoG5Lqr5PBFiZX514HuG2XjYe4JsCUImkAJXXa1emklIoILycvS4hN6F1g8lwyCle1Hp4W/eG
9bJYd8Y+YyJznWzfmDasCoznK54U64S1z3CQeKguTOVUi8kOgFX8xzxezEeuXarYhYU3hazQxygi
kAv5TciYX4N1Sw6UWjGEih7yPQyHRM5UbqiY3/LTMJ9Ic1eLXCkOCQnTEkOYdaF/81BbEwCQqmro
AuFqZav1mcKq5ZJDqpwNmk0FsqoG6aYWSbLGDmxrpeBN0RrApWZC2THFQX/BXS2vU7ouI1Zq+crt
fTUII8H046+VoW5rjRhIimyO8DAyL7FKsT7MEmveHCIxW5vv9DwBBQVwq/ADS4dQYBcbyr/pkXxW
xTxOs+uybIIlEXf4W1paLfivoeWwoUHb9skkbZfJK5Mdo4TY93o1MS/18jKV+iCvG76h66VL6jV9
7D4pQDt88oXxdT6nNZwouHIcXW29hSdUA0tI6boUeNEpS1FxW5/8qZrN4XN991NSpSv21ml1NL1y
Uru9zx6ZKsPky0XvnOQtN8Apghrb6lNMLQplbESN/UxwI5Ozd+RMLINE1x2Jv7PeibQqE85rAysl
HRaXw6X/I+3CHU3mPFuyoOEVkN4bkq2Kirmi8aXIQG5ullY/8ZSXrbwbkklNoPFqE9Gx7WHex0re
HqLxG+W+X+HmauzIZXoBDhGsz8JNvDubXoW20v6wVnVf3Vq7CQK9XAIZDJZv3HqFwn1YRQS0p0DV
QFlPztFM6hgR8ebmtQKXXF+TNZxjdVlUb73TTHIcGt+1yYuj3xV6vSUFL3x5uFBEKSt9oJpGCyGK
UBd3ufRDMrfx36Z1WML+NXhCBP3vR4XHN7tugednGKCnrl/hjnJDpvqtyfZWA6wywkKSsYGeTA+5
L0S7zmdO5m3AE/gjjL5Vx3LHzu6C5Jyj5wvMTQzAvNLaDNroT5gYrrbgPhKxjLLb4VcQCVtgfgJ+
BeT2sRMXWJ+h7C3SLiRPjmrBKkaLshDnAGt3wVSSMrEUoQHoze8/89r13O3MoDiVpxWHoX74Imej
0x1Xg/aIg3Qp2s+NjJY5gfuOa/UMBMpLCUI+kESLtCisOPJY0RSw8WXSuWdj91LgEOQB/mah5INB
vj6SShBCiB7PoVgdSO9DVj7KOoIHYCCxSLRfMPPEaw3kQm25OqL3YLKz5SeYi0ZHZs/ysje8vxH2
uz15ezAazOHkOzkXPv7ndBbUgXYOv4wtNx4KMfnPD2/zKKHDnvUQVbbEPB0H+MkEUwgPC0h9DmYN
OVcroF5VGEj/TxGQcD0ujnxIjsJ2zNqLGEiJZSgpupjpTUxEu2aYpySxV1QaggnbOj6iVF6NBrV7
ObPCJvs+1tasFryPDzg4YJ0Z5Ml2EAB7cqFt70hu+CkUudSmbn+TUAgTpuNYZ9wz2eV3nTlOdx5V
o0rCjkweP2Tkn9eW+mba+pqYqJxr7qcDBZg7g4Y4kMZwYr26+6ZRN07rSY3fd/hKGsXpJ4GpRMRM
JGgI2N+w9BsfQw8pgffwuVZ4MV6TdqPTSCPXx3Nuj4f2j5dZuoJU6fmjHhWm5SZnj5LiNDFohLOh
FGCXVDBfJnlU46bIUaYljSzzA9/yYCq90jPGzOJJ0eueNo8oOlpmNAjaHkKUbxmOuIker0XJFhxR
oSI3FDFVwvMMnjGRjjRI2KBF8jhrOC4XyH4cpfn40F3YQo4Y4tb2CVHTCi26x0jAW7BWv1lx66su
xdB26KDoi6uDtDfqEDYYGgv98baKS63byeNPMLGyUCn5CgPsP4qQ6AxPJUiI4JH1T+8j7Q+d1w65
wcotpx0CubYhsgch3AWNMa/vh0dk0GEA5Uiev4hyYcXdZRxwI544H1Sn1JChZ37L8ma6h6erEVYa
Opr2iPZN3ejGXPpsHdQawzSbriJ2RqEmDbbLuakHCueTT+6/+V68sO34mA3KA6VDFd/7fuLKU09P
CkNRAg33B3aqSwgEfJnQswq8PW32Jk0AHGr++0bqdVBuXvRNIKIXu/kEWWxFCb/ItONceIW2+xaW
wiShcx3oDF49XIw8QStwUegbIswMfKQIDUSgtIEJDRJeQy2rtgAErxz4XGJ9Vwyd/W9WPOeBwoSE
xcdHb9Obvqce4MrRRKvP+QclwiYry/Zv1BtKLVyd5r8ahNpezHEvahdb67u0n+pnpWsJgOF+AwOu
0PJ2zTjrzZUD8IRsLmwKmRWNNkks4dN8OmnuBB3Tn/JKMIjgKRM5hQDyCpuWIWJHgoFnUiV7ayWU
xH8VoahyNPs4HRY9P70DjhOMyjATaOATHm8p2xjDpUpDslvleCrsHu9V4WZmWe83y12zM+BoY3HO
zVH4UfBdcJ+9wQYfkKXEOfjMespalAvHVeS4qPSn5HOCCvHK4rmzIpvVBdWiQ4UUo1QtiKTDs8xg
n9mRy8GZFwy5hNEZWaHU/r7qTpMyx6sfPJJePlazlZunDaZOzlqydG9IGwtqT9VAidzlW6gElDEL
RybEhKQac9oAEL9nVHTJBARI6peQ8fm4jopPP+9BQ0VV25sy1SrgKkoGpIsaxHEii4qHYWVh6Wsc
K7Fy+ZB/Ct9anjYPKWr0133PhPhippXcuvGIkv89vmSvR24q4BjiE5kxNa2EOyhzp36CzZXxcvi3
hpE7r2fl4VSv81uH8WojJw8z1HqZcbMy10//h0Y19WQpk/5Erovn7ugpJNaVkkB21xu9r3vTZhjw
2y3cNCa9Wbyx3XJi2L7x3FoX+zrt7S0nrR/xJ5ytTdbBxrEKdgIeZQl9OEPblLa+XvTVKwv323Z4
37dW4lU7lGgN3Nksf6t4+pp+WeEdShJZgqJFbXq8gHBkzLHM7MJIuK2QhMX8THRDL2FAEHeo6s6o
DNveQ/frKOftfe1IGflW/tmeK8YG2KGr6w9jzEhZNymFcorGlMniIPbBgUsfcPuQYG1mZ/db8K5L
tuhCg67aZWyLVHcb2CGxc3JbQWGLurPbp1Ox4zT6JZvf4YbYOJ0GS8ft+BPaqXwXYbV1aTilfzma
5QX+n/V64fDJP2PUFpdfSU3uEpD5/biYoWa8r6O39SprV9rSbeRBD1F/TrmwXmL6KJQsfyMDPZL0
4deCHMNw2Nwig+3shF4F/fiPtfIwzUFfWdi03IGgasL1ZpB5X3UnCd5C/YV4k35YG8/KerKhz+0j
J+YqePZk6+jFYaChkVF9zlnKZFpUUGBXEd058JFu5groae7UxFz+dkF+2iJ87PEkkTEGK4phjk9m
ZE5F7l/1Ai5pjNwOZe9rNOfu4OgBGSQsQRQ6TlcseH7iliV47eDBtcVoIQ63cLGrnxuqmVWcWbpV
fXZT5IMYoDnqw5Op+7G+aoUZV1whsX3/zz5dIIRnz1erVerY/GcgrY0cTftWe/K9Akv+ogJo7A8p
tXI7RDhgF5FwSI3t7irbvA7gI+696O3E9MtYk37+53OsM5TUOpYiivH9aJCCLkeP0bs0nApygkyx
2Pl1SmLAM9Nd3QrIcsQS5ADZ+MgWCTeNmzMtxxjBmWTFYREBXmhMj7rqqWTG7DSHVWLjpFPuiZa8
T6PwnD4rumArvFiX9RMzGU8E6v431BeUUhlU8NxEy2dtoQ/2kHYUKzROjMrt696poq+gmE5mzIqI
zrDZFCf1Fh95KV0zzSOury4sv4eWfAdlXkwo2YnYtDJLclZT9q0+DPOiKRPYOx6wi8j+FAQR7dYn
H8Wo8PpxYgnssSIOErwPyAZEjbWVcacfX1J0GXsC8+phMiolQ+4hJgNQ/UADXqcgRFLIYg6p+RXG
pXvfz2+gwHNHARwybpOZzidTRnq6gwRNlx/SQYuSFKhbLO0huSuFkpp48cfHibWBenEaZdUviwyM
QtjZK8HchgMPEo5OyyHRFSeFN6xUW1BVQWEJhEKIXfA+9bi5PqijOYvEOT+xkahqfwxmcJKNWWS/
yyG4eLnioMJFpmHbvUcA6bGZXd6268ZJyKXkO8NGo0OQmTgQElAJrGAPmJ0GViNZQ10NYeiFJ6Ty
iTr5yyr9I6MI9+d42MBwuhWzjZ2oZCbqgmV62ctpyjHvCy8fbJhBVlODBjFiErtOZRixDv7LSh/0
Fgp3v+bEk+BNj0v361y/FXv7n2Yc8ibQzHM/c/fNyOk+4FsRk+LdD4SGOSHQ5qzzd73TEjdDkxEz
ByJFJ1dk1lDxI76JaqpqU2ZtyX+OJMGUEvD4G6YoDsJ4KGak8oE0VjMs/uFBRz1OM8L4qb5lzTo5
WhTNHnI4SficEh1Mg68b4/U/VUJN+uNaq7Y/kT379JVS9nyDbCNRBatCE/diOdZ5K64qMD30QrUc
WdOxzb4Q6ABpWIF+RKIxE5BRl8ntfa9nGsWMDGqJDKmRvuRBIitIAmUNbe0CVuRBG4A7akCWtDcv
XA4FfBUTOoZpEWGHbChlpfT+V64A74v3UlDnqr6u+mEgF+UvBW+qAvxrTSUrh/DYzXjTQ0Xcp/eo
kIhit/SLYwUEQSLZwIT1LIM/MMzSqnpQDSOjdO0DAxRbvKRAc2ml6x5L6/pynTnipOOH60gxpAwb
o9QYid9kR4QQxycKZKm2JyE18j8o+1Op3K3I6cnw2haczAIEK6IaOY0C3ElCcilWzrslyAeg7QVZ
nso0b3C5UpOD2GFeq9yT6DsdDZw/gOaQhg8r9AeLxlcPUHllfI0jreczkLjQzCWOkG4Z8B9yvQyi
aQov4Fw2gmLIvl76uS8Gw1zxGKB33QTo4Jm7Gd6jXxR0m3r+/kZEdeunmFMOrXxccq32pvfXKx+j
q1ptFWO+4YDHK7hibw1gAgAd68Od3QPkvyeRrAl4AcFyrlN2WNuboakTIxCdgKXKYTE9gKXwi64T
zfp3uFqZUzG4iwhkAO9Xb7dUEOtAqiv7o297ObUfs/DwhC/aNCCQPsE5j5maYoYVoo2On+0s3Cm7
HCcx8fl8yafijASM3zr12NQxGf6yq2F4k+3mVmxOyftdCJlZFpnbMw5C5OcDHWCQ8IfsNEMz+Bgb
6sBpm1CZbyZvZS8JzqTxbwbGFGPZc/D8ZV2Fzgy9XwGkIqWB+/Duz37t5BjhpF0MoW5Tr/WLf9B6
8MdSbtpV+p84ksmMAwlCNeMHF0CWiybv9HSuoRS6BfTeuP+25/J1EF/0UT5JNpD4Rf0WpbO62RXB
YJtqrnf3XaoheOjiGjk3+s7sn/ajMwu8IKf4vXxn6UyRZhEQbh3ccRvtG88jDYA8Hl6OSDQwFO/f
nNhEw4Bt2Kbs0sxzzZmLw+h4ciwUWs0b6bfg8sJByLdEbkd6NMJcdL+HSM3iQt47itfbHRaIUlOw
kBcBDJoaEaa8Ke2nWA5XU1WZqzhUT2/VEmDQ7FPYG2vQ1cidCYRpKWrHDzlzIKnDjQIU6wAmydJq
bYDNhcqkMo/rFbRB9+wb0T/aZbrGkNvyYw5YymJAflRkQ6/P2Ru+qFKGWkhjscWIwkSEN7YwQErg
7iv7EzYpTzs/sWzm1NSIdAl9yjSw1iRx8E71OBdK4EmKW75T1kMCnGWLxdGF/alwTEF4tJWu+uW/
59e9xS6ME1oeFazMBO9cON3TU0hLQDqMuD7zuBsERipcHH5oJ/y9l4pf2W8FiPzrtX6EUI/KbpJd
LFQQeb9Ujm5UGDCBQlv/FU2w/EjVw/SaSfUHTPjLncbhKkIpCHzUgxP7/GGL52R4eL3nl8iop/vc
XWjj/qmXNWozJgUe1LvEWoztjr7fESM1GfC+ooYNaEbseuuWTrkuT6mOaSCNKcRsqaG+hlCDRwf4
pdOjig8TTMxbSTrqKyWS/cBiwa32EujIuxJdNS8Ks00jGiQ6EIucEQ4NkSqMgV+iVYClh/qudrE+
JgCmc1YvK5h7AdOeS/AXO6crMZadIKIiHq5+RQVK9MQLTlTgGJr+FtGnJeWkC/NY/xX3uYRcMYPA
DddeU5CaSv800orGjpH7/bAAl/ejIwWQpXccLYBHkG/PUp6aLDWyBZSTc18cAwnA+QkBHCDHzF/7
IUWHm9ARDOXcbhSZZeIismNQUyZsze8JYFnKVvUEm+0xgzNUwDtAQG/JkrJ94nBc++Cgw8zhWqrr
cw2j0i0NtDsN72RflDm8NpjRgv/1D3dlAG0tVzVJmR4IMPhPRlX1n/f6GMmnSIkXWhAkD1NKS2dG
zR6b4PR+CkDYr6a7z3ET3/PMk1MNl7WLqS4BAceSALlMpnXTLQUIG8OTMdBMlkN6BxbQoOosaQYo
nCQYm+UAvqs6LzX3h+9GJOR8MyxTT32HU7+25EpsQN9D3tkC5lXvl12/NMr0MRJyxgdqCJUGuGB1
NlWcpsk8yiF4AUtmvn1UnWyPBKRKlBwSps8JB0mXVlI1wx7W5JVMsk8v5+CqLfdojwTU29SVHMYP
aCXUQrUveyp8KJtItAXgGN796JmEAUI+h/XLQayM0OSmiH5jT4OwUjzLoIZ/P8wePbqnZOxZib2x
HKnlK8DwucTYQkqQO3MCdiH9BN3yhAowxzIE2uEsFDOXsZgfS2CKAfKuKeB1rxJ3yYw9nCTF3Y0t
KQZEFcM1PMjFZ8ww0JVIuZLniTITj2pZJB/oT3xLrYD+aUp8BxwpOqQRR10NEB41m0Fo0bAzReEb
D6vah44ke34fsZnQY62fblPa5pS8Nfqqcts57XDDN81JH3ZsABnXbd7SUANpRt64Wa32y/L55zKx
E3EToP2vfKfgF2G8rrmTSk1Wbk0+vnqymqlf2yALecC/bBjzjVcqted+4akDWHzEozN7iqzaXr+X
jHKTbj77Na6gokc+Kdk1feUWUCrgOYjZn9NihVaXOTkblhDC6F8GmZN1wKDo11GCMcakXd6IUXcp
p2IE3iGQ44ATQ7HS9kiNES3Ou19RLZpdsbBX0yn96Sq43TUpo87foDEd1SWIL0lITPjmvyB3s5kO
IMUSLIpZU2k60/yudzQSaEShwZ3ydNQ/okSMg+evSD1oO+F9cAp7e9WizQ52fulRcn8bYIueFB9I
UFFvWJzLmPIVznVqPtKMRPfRr2khFuOAKG0n9Twg4qvuZBoPcyttQmJe3HpAirs6qm1mTaQVSXtM
USJ/dMefTzB6rDxcCaQr6gjBZYns4ve1VcHbT/hZFFvHZyNJyLgfVTZwP15U57kgCjUpgzdTR2Gj
sb+l61iX2fKzg+UHFe23URvLVz8OX3TLwvqvpDSKdHuHB4QE91yKVpSJfdCuEFCozm/AABUHGLHD
gWK23FC1XmBTWqCESmOFDZUUuBkUn+pdDVYs2hGoTOf9u/fhd/S4TyED6LX5FZoMumZ0K/T2/8Bs
uWG1dta3Wr/mrDAdNFiSfcp37jYwiMPVx3UjQiZC3807fmO97Y9ooj5iwKZmyt+Y4cP5kl8ucDW2
RtlvZIOI2R6UgPJrQ/LR7/ysbC4sA2Ig3QW1BfUaN0BwUtB0YIKu0KtSp01ft/wes7WHa/8l9okR
Psbqaq1ZJ59htyrhgZ17HzvCBUs8lvH38+GLN6fFwCsxJH8poRYFEuHVk7aBTu6p084XD7lqVR7l
MPm4ZBV5Xl0WcuV3qvqsnWQsl5FcI4EDaNcumx5OWamuHcW77sPXeXHIwu2pCpLeGFQtlNCl9sZY
pVAE/XrN8ua4cuQishfG3OahkXiiXnjxo0Glawp75ioN5QFnvNZAiWAL7jqyY+f8ZbcHBUjNd1tZ
Bf5pt33vFPXb9ugNfspfWjaE6rntEdN5yVFy3JgzMlExSUjv2Zfgg96GXDkHzs3QrdoUflP+yhfP
VUXQKqi6rcRYIiqjPVJOv5tAbZ6Jz1v3p5Xy5gZvgvIJjl2tGmrnTSnIZC2fVWwkIaM4apR8KJR9
oSt93hR9GidNiqAVEp8lo4A6+3STtrUhVGXbghvcRed9sjpewhuZ09A/qQ7Au+46zVn3QXLdfZe7
/kyM9Lt4jdWda0IDFg/qD/l/hdEahyynTm/HX5Rte7KAx12l2IjhgZ6F7n4wVGHVRTvgV9fP+JmN
6jY9sM2SJaKdu9+61Yh79L13sCKLvJ1xickvvNH9XL49IHbgT76r7ygpgDK8iuETx5rqizu9+GiZ
v4Tlk4gvYekS04M2ps7q6kbo2A3WQ35aTQ6Ssv0vWpzC9GkZd/+BWnp/u+JC5PjeqHPyyxkfnobr
GIRwqFY76aXycCTAKgHCQFn4MqXN1DRbo7YwV0cxrbxkpwGa9d8k3ReBDpI/Rx/UshTFoEaqEgfa
4ZPw0RSiHwtxcisj146TxPtkNCkMNGGgkBsvNYbqQ/upVNqIX2usC/GKjmr8Ka1XZvW+S+PA/GFW
Ip2fE8fIKdpCd/n3Xi6aV7EvJnsBpBQQqXLzOOJOQO3wddC7eHhIHbtBryYKTwaB/8kPFwwJcgjX
OYWCpvwXacvBrgFcs09l+7l7IqRNA7QsZQFVZVkYsyWBX3/MB0eOIrzzFdYPnGxb90/E10TPltcl
NOkEfPkGy9PoF9ak0+06uzKYsIWkPGk5ulZZA7dDmPVRj/rQrNOEqX20VNbgsdI50FFmsxSUFUQC
e/Z5fazyeL1VuTR2rQoblxebZmrrK6UQ8TE84SfvV+UPT69ZSX2ZedypOfBDVYkyVlhK0ErmlWW6
D4ENDBtJg+ER7liazm2J9g428fDEIkhZzIBoZXKgdrLUFmZFvccpKAvvQfhmaSvZ9zihTR1TNuz6
oerDSFxNen5sRuPZzN58M2ySWRxNgJjzwWC96gXNPaeTQR8usZ5y1tr0hTJC8pZPm1eLYrAXnOlr
ZIHKaxIv+fUkXeq+J9NLHkHpgJjHp13dN18GEfsgrbg5xKVc6ZfnVQgWZH4W+QK/jskqq0VwukxC
utFs3+MBxAQMjfD1hW/6eXVQMjeAZ8ucgaPMcW1c1IcQbggLMyVKJDOnPDSCmj+3q4pCsc3JCvie
6rY3X3pozXGEk4SEUGLsN4dH66tLJtbXLIS5BVgJ7bSb+1kak+5InImtta+QG3tuVd04CXxFl5sm
6FJfit6G0zKVlq6Cuyg7tHxBndclaSA+Z52ya5dR0SqHesQTqXt0+xhOe0M7QA7SAMTiFuG5fT5P
J/LFsK4HBonJDru8VXnEuaiWvlF24IRB3VchCqDY0Bph4VTL3Lyta6rsOjnGRwizGiXREjs5f09g
CSNSTPMslv6vyVeYcuMh/axq8KqqvI9gZTTWFNGHw/pobMVYI1/cTHCualHzGcZtNxF4zhmLpOCc
OO4X3Vj52YUD69gQ7FyxaYU++DHPd6u2uLGzKXfzHOKv9izRK3MtFdi0Q/rDw9r44LdnS69MUHlZ
OFqh0YvqRO2abncbm5frAWvcMLuWkLIGMfOEyZnx9lBvBvzSYgxs9v1jsXfenZU4ft9QRUj6xGBu
VaRdhzlztNldem8I+AiE1dZ9rNXagMZvqGHCHOO2tbyRPQbT83ikRz3VB3S6Dl5psqFOCNN/a+T5
+55W+LsNONY95xBhii2STgRFkTmBTYUs3xcA3BYaY8QbC+Pn42HAg4x0Di5+ErWxCsZYB7vykG03
y04hkcVZLqOmF5b303ZjLiXO1NgA/8m+lcNxVA3LAc9UNlQ6oxWTcVv+5bMAUGUx9UXFPLsoCJyI
9a20+dNxjakRxyMI7qvRdAXT/luSEqCJpy49axsIe1hyo5mETTHgFaUQEhkdofnYyE5+Wp79/4BK
wo3e2mEbSla1nj2H023Fgu8V533zyXYdO+g1Ix7YPk2ftu5IaKny5SHWGf4S7OtVylRpVO2tN/fM
TJuqPcX+9SX4ZyMmKP0YZnHZNWwSDKHm3NF1/WMBDxh5S/cimv2qcxTmyt2uv2UuHMebNAXUAfKu
Qd7rGWkntnlWRFHIhGd7o6ktSs5UzqJCiym5Bwl3tXvR6BQ1Pv7CvskJEaTBSRI2NPOvG/5XxIJI
U5MKC6nNqCXTEVcfQTGaMdLNKNDLxJEQaOsOy8uMtnC9Gldg0pMnj6bm0SqE6mjPGbsMqXPoylO2
xl4G/YSIk96xKdNk0ZOoYhMccO3tHu6yC1RVfHeC9+jz1NvFCfb2P8pxVQKClxxJPoZzXkQRNW0T
vW7iw6mVARAyjLfOp0DIWf5hL4gBa7ImVhcb1hpTPGkWpoTwtyDtbviQL6fiadDGnRZPtD1dH+Gy
ZnNQ9G5AomPyH/02ieiieYWDv7xH/vp8WKfaLStfJ5KV0Gcc3lIUItP6olYGdm2FgIa6H2JVHlTL
COdHpQWi5MTeSoWt+bKoRlN7PaJ+sduPaDt0L4pA5XwkMGw0fYaISMfi+A/CCuq1/G98uuXZu6jO
KghGexrgi+D+XCOf4UL+kTOsDWD7vqWqSuGw4eoq1e90rZkAkfPPapst2PTFogfING91F9kCI+08
r2/7qi2dwtd6Ni5rbFnec9fFmlXAWr2ORvRJ3X0GiBX9XjtBoFK1c9JnTX/fzTl+p5kDNbRPVMW+
AZjqY8nKnn5Nubaj3GqAp6e7GmjxC06a3Wj+MaTZEgh8fR6rRBo7+ahhgwz5RN19wTyN3p3zbfwT
hRMrOO0Avn1HotibcieBBUY8uSU+nJ1bnarokdMtJqxjeBFlGYdT4lbuKgYpD8iZQsTiT1NmXwHH
KQFjAmyzBs6NOP6P73VUh4+yAEQCSQX886l7Dujb14w3fXDs4RSO0yio0KyYOE+6gQCkOPYozXt0
fIvi8X8feUsCAq0uzcgxWbANLdGX8xJuT1LheKdkxsJTq+5iRYq5zWho/t4bxpGe5PANjnZIkEQe
B3v1Psu0IGfcqeLnoahCj7vJkOi1qfo9OJLwX3bBnQqhTQ1aXieNHQ17fw8tfYeuIa17Exn2PGSo
vZC70Wn3FL6d4ErTn3dQEOR75+pC0W0q9OqvDFnPePGG9JInLYdzy3MKDFKm2pLe2jWbnI0KG+wQ
6Hin2/O4au1dOSnKEnoyBMBubtiOs77nhJikxZe8Cj0esvJ2Ee1NpKWMQEABRuDeP45k+RryJxa4
SuJdatqRAsXcmnfy8xYUR4R94qFv6D3BhtDNMS/nlz3gzmGjf3tSEb3fSjP4zFj9Oe/nIodKt75y
lzr4lCxvUoSeomqSHvLevNg9baao90c7C9xzffNt4E7YR6mZHXa9Qwh/EadXFvlNtQFl/qSMKk6d
E1s4voM6S+FMnV6x95k7zTwLq1xsWuDn8YmWyTyoqqx39tsvGN362VZLx5oDynZZOnuz5e0nT1ZS
jS6xwvmtbWZjIwqTl6IxxfuaF4dVL05C+ktU8/ozRfcYzdMWipv+4610I9DOXqvBRUdJgeJoAiGl
oAhVqpmk4ShJLHHBw0gC2IBMr+9KLCeBdeFhPMo0gO7tzkz7Prnpsbdje/Iz+/6cqGuM/AT3DwA6
3lU7tVMs9R9AG8PxSIxaZvtw6cGsG2BmUOSsgfOtRpuzLZmFxxNDIcr+T0mWkoC0kt4YFaQnNGFn
lHeR66X1UH++wXN3arib2RpBm9nAjNzP5EkFTFgDkXGBkHy6ICm/37sExKXfqGQjCCKd7gNKrfhp
oUtYP03B3Tf09nFVy69Ad8ETai6AedEev24xi/bYvIJoMCByofFNZrUr097c8eJt/uofYvvnzDIg
PPFpD70Aj0X5kLsVIUptg7WWw9G+FFo46x9RLzNqH/AtGR6Hy0EAWGAhsM55wSD35SZudr7deE7x
yo8C9S47uynGH3a6RoE/MVLvkCI1AytzOVpSjg98v61x5vxHCAhD39HH3e+WEmw1NhLCJZCu1UYA
FyPQhRMwJBFmv9DguRcO52E773aNMPqam3szg9A4gavWT4Jw5T2102SbCxa1SFntayUGugG/pqGA
fxqRgOzEOVJA4UTQa1A4HHTCHbWmJ05KOzncAlssIAHEU2G1gESd8gpKjbIseqxCsL8oUBC3uCzR
u36Z5mDT0nT2p+Z6grfSBWO/UZTP6jGgd1E6NJUj/ItYV3Kzw0ZzCDuhyUCaBAK80B8VlQDWK9UO
DFyC8o1NuCswjmhwrOPkReqZBDlhqUoKv2vj48qReZWhWZdNc/+Uc88LYWiRF4r3IC4+5qIQ+uLm
yk+OGoJ01F7XS38pLuhIE1/6MJTrMvSsHZOmjoITomoc0/et/qR8RQQznt63GAoK1fwIrnGucKJw
he9blMJJEJLKld3qHCVCvrdmojs40iVlkaScFNBBinymouxPH0QkcJlv52SGvfOsED8K710Pow9R
VJRpTB3hZFNlBjStIebqeGXme5F91hSqbRLoMlKvkuo2PmI4xImqhR7EDI6kE7p/dZIezWWdlCNZ
2/qqMlgqNgme/rttgH+StAydZgYTkKKtdDR7wVXNu9D45cxGJGLzXbPxMfeMwtGIVirZyPDwogFm
mAocfIkEwcYL45Ds8vaFGneOQSXKerxVy9AAnHn+YLeoZjAvMedt++S6/nYi+6Z5Cj0aUiuAya6u
/1R4cTGJKTPPbOdhearP2vSTCSxuK4Bp1Ep+0YktV+6cV6zKwFYmoQbVtQXGk2tptaKP+fwFzbAL
zE69r6oTqR6vFgiDPBbOipfpwjEAZJvsh1YbkrtvmaAAKstgbyp7wvmy3VWtMx4g7wVYAls0YbYS
8K/TKhzicm1QO9lQ7+5gMY916Bn7c4qTYnKBHKJPq7LNjGoHoL1SSR6wHwMvwKvoxhrd/smZV0bx
C3MIIlGfPdT+rpulFPO90w3SESvkZkSq/8eDbK7gxpYZw2fqSKHn/vti1oJBsgG0wuGNEZglCL8L
M0+32YblA1RxjeVSvsl/q2OTWJT/C+DUXBR1IHg9Se+Ofk6tEGlTBSbKJM+a7umdo1wQqO61Pmh2
RWa9/zJ8a6bVPxFBdLwNmX/ziXu9JnjAtU80sVbaPgb6PKTxX22Bly1g3d5ApUm8qG+z9PjAjNxq
pU58ktJBHds2DWWSqxGAhc6qevelwR8THq7Xzcd4IayQFbUXsnH/UhqgZ1r6JdusoRr8SRkXAjis
gv1KdtOaUFD5IhuddrBkqGG3n2Sn+wm4/1SaUw92+QtjY1sVUOlgVhr3MMe+Tcgu20OfXkG4j4R5
Hz3Cq7d/TmJxEEtMZiMJKJ4fyiiVS9OFPN6bgCYK8aZcnrRdoD/UNKTwDPHsMYWH/M5JD+XUeuc5
DB2rcBTskB0gXUj0Ny6A3dlpITM9mYlb3yzwJ//9PgMd2+p5Vh18B4R9l/1If83WD6/eK6nRdzNz
h9hOYp2NAmn7vBBVrkumc4J3PpTcihYImuKwpV+821EfiFSob4KxTq3Y/ItIbvY9tjxrgLdb+Vd9
0qeCjf9h3XJDjdvh5pPg5tEWRewqLg2MeFOs5V04YoTdUdhV4bl+dCHxVKvpXlTPNpLs0CKHlO3W
O9nU3fuzWPRRuiEe6u/o2EATLOJ9lPOPB6xH3nE3r5wEWg0mn2F1rUmdkpN2fDGv4z3EwrQdCx64
TnrhlrUAzVLjW7E/xaY3DjNRTaTDagk9GBrUbQ/F1hthiT9EKU/Imj0Xb0gISyO+xnMqvQtg9VP0
D63vdo/HtK5GryCUI+AKok0TWe0OzfDiuT/ou5CihHKdsKHlBJYVbLigM3NloYsVHOLut2MiuD/v
B3OdVYvWtoSfLFQYuzuvtj5PmcNXlDsaLZSsto+vOCG5dBh0uzsTADZ00DMxNMWI8L+Vdcd2WekH
fQDCTlJhoEQ4ehNxElmm78PFmmecZL3xnz57QK7APgcxfzn/Z2ts0D294zgHwoYSl8JSrTABcxsd
q9w3mR6+TwX6grEzn0t5j/wl6DtQiWnvJiEpLW4mpoQrT9JqZ83lHWylGZFrpIfjHKeDyER4paIe
FnWB4s3mCgZoR0L2ULHtqdmCrVWQJzyTuar5VGr/yRUFSDUhrOs3ir7Yqj4bexEbQCs139mYqhF+
FQHdOZ0wE76BRVFGDzfgNq+mjVAhXGORUAbFWUFs6sjfXfTmxuNS88JqB7R+EoXOAX4rcqa41chw
wsKEdY7ee/d74p6DSxIr2zjEwe8FrXq5U4JfsHrcTgnV24ON9ElHKv8Bz1qCKz3rOr+d10SK5bFf
L5QixcqxhqqhriPv/i72eG2fOxPhTx3e8/xrIfDVE9sZMlSI/tnlnJ/FLlsVz7WCMUvRCQT59ogP
RBDE1pyzL5u4D2KVVddLu7p7JowgY6XtBtEzqnQ1d5qEUZY6G/EkxBoy/rrDrcGohaO0Id/SRZC5
nMSe56ffHP14VXv8RlOV/oFYv76/NQdsXe7xx0c9IA2dVGLTOftDQ3SiVopfaLq5zhvHauKBddCO
M5k9y2G4ItJ7hy8FPBdidNant4YEh6QmrLQhk4iCRXgvW3rRqfuh0lbKWmugnY3rS4UiBslMBBve
Jp6daVbMMeqJG+9OXH20fir+ub9xX9gGMBJTZjrDIKWjik4hCAELwAAzMvtD1qnUEHPV1xk4nvJq
K+Q07f9DhIpQOVSQf+3j+HORs6Ye0Am6HpFcqmdbCtPw3f8S2IZFDbUGFfI+w+LLAH3sHhWNJap4
xhzsGyuv/kjiNDsW0TgdNN5uddJRYl4dgaLy5LkpeHnXF6gtp6jbiFi/feQqULa3Jb5LsAbyGbcx
Nfr4XMlZVhA1fWSlmmEeUyY8K1p/0W8LFB5F84KAEA7ZvRE+zoR4sGF2qZcKlljWTccPx6X9eiZi
JUQjj7mJCf9KL83SlASTSNYOgUKX1Yh1PeCOsERqDNSSoTnbLqozcpf+8wvFxuEtHtNWqqoLmVdT
43DYjYCLKIIbZYL16GWHMWlMWaLxzESlbS199rD6OvCaoPegFgraLjMMSt0zQi2nA7mlfYRCNUtB
6vmLtBXxRk5M/28CfP9HyrtgqhDuxvUpaWj05Pq6voRA2L4a1vMHK2f2b0eYFRhRBaeUzZzD05qe
tbXacOxTK9ZiP7xeCSLhksDRJIYDjQ7TZnqm7uLhCDE6/OpvTwgCZ+bG42jShhaqmF/xg2uvCgNQ
xBS7CDPvrr1W+PzeVq2DsXMZm8ejVBJrS0heVwo3cgUZTT6MOSZvpxHXlXvBLY86CyUe0jdnusnu
6askX4200XoLrkjKaTGcTfQ6D8tOqEXJIqICGLgX9ZHbbTIoNL3onSoLKUZODYgL1A/dWQDjpB3F
E8RdCKHL8rm9X32Troub68Pkr4hBnuR7V3Jf116N0lRLME5dklFUcYXW7HinVIpSuow1tl4S1sfg
bTH/Z4im12OxJNmpMlhWwBmQ75oqoI7tCUkSmfPztBxDyWXqMKdAYQqajXV0QLjO+u2t5dtR60Sp
SHOuu+897YrAnRCnxFs/7iLyoFaMC6+UmvZyYqkWmmNmJuofUW2Q7WAw+7BbIuLxDWS+f5duNsav
7VI8U5BbonpiTkc8MDdVRkgs91IJyQR5UDuVCWCNpy2zTk8JIjzIbYI/K+LXyAgf+PQVxKNg8skv
25O26ShiyzTACJPOIS1KtXjS4mPbzCCkprkpSx7bHkGMqbmhBpIHli4bkz9UJJeCL1yfdKPlZf+F
2d1bTcI6+/tVXtHtvhX89RALgPeVoX5DZ6SGLIZU+iZnInMMADSape0r9ZlZ/qIfFyW3pzSfEedT
OJAYrG+NvfcSGyE0J/1qaU3dqt+GYGkdqi6jrphYj1G4iXwt/vTCUrtS4b3Lhtpy9BIvEGdXEJ+Q
ymndTkNkHUpj18y2UT/CXNqQmHBj7eBpgTJakvxIolQKTiNGrj/5+cdCBZWwpeBRDlLjXqTR6TJ4
7eezcpH9r6fHgCe1lFeoQoZ5BWvMvcyrVtRf1PzMrR/Gm8QRPXCJefMEnF5YBPC/l/hEwAg5fvSc
mmiAk6kyKNUm7gRLFUO/ZPtZ0rugmZEld4weWiz+NFCtCo4X1txDlLUgY4Ww/DWyB+lt+0iqtEU7
/aQs28ZZjg6kyGtJfn2weEQKPpwbxTXa8i8WVd7ojxE21Rx3La+ARFvM707idF10WfuXlfpkSBYR
8q7ijX+MEKL1u49hwhJIuLlUgNZsBcom2Y46An+x4X2b7ms4cfJp/+cru+DdIiSfuK9OfGgoBX7G
HVYcJcSbuf8na2EeMkIVcLCbEkyUuoY0Od006gAl3TGpJ0pODlNFc4dO1JbtBUVpTr00RiAH6tHP
WPP32B+4Xzgl1/YI15XwIp6CaFGBbovYhTAmoeCzAWox+e7akCHcXAkfSJUxc+QMaOmz5C4lgrPV
mCCJx9iDJmGxJjePqc/IAGBv6P6gMZwf9YnAMG/lQQwf9GSri6xDjp8LdeGZjR5+EK7SOu8jTH8o
FXpmLD5VejgoUtPVeigREofe82yK+wun96Ld2/LypPXZ1QCDfVztOIeJP2aCNgHvam1Adw2Nvz81
tJI0TrkNClU6ZtPwoJKkL6EzkMH0nXSlrYfLb21tCkNfeGomVWPVrGNE4kdOUFKVQ5TZ1VpzOlwZ
u/lSHzNDTy6yD61muDy0v4/EIejzh403FcqTh/OvDQ86Q5a7KxpKYDVJfG75N8HsyDL45xwbs3Hx
V8pfS3/nfGjb5KdbNBD1XEm5tMV181bP6OpAGU6OgzFDbHci6b1BcZV4nphGFcE0fc9bdTYGarlh
MeWBVZkprLnQoQimcndWhOOU5Q01Ul7BO3DAZ/sx8Fm1/+yYzS3i/nFkaWWBsi4PXNvJRQtVsOsQ
g1utzF4ih4x/XlhqKBWQQjp+7rIRkZlmQltc1UjTmhbj9hKjJxER4Ka81oFN9pXonkwapqXbYqmc
zNa9Xf+GHyZ5uvAnib7FY2N5tDuiTfRLoNbVH3mvRFUk0eOB4sZLu6lDi2vLteCozz6VgcWTyH6k
IZGF99qz4Rzl8R0XnbLPsG0Zm3gkkF+a8BEL7GxxlafoTj3x+iWJsnB+dRBsWlaDzKYmk+MPJIJN
Owa6y71g9oLMCY5gq6pjSf8pTji2f9hHPehXT4CQk3xWfGGl7Kz51/tp5z2MqI19IOyfL16nu8e6
cRILXn7JlU9Mt7D+gyJgYEFr2l3MluBVIH4Yon07wEL3EXox5Z60CHVPQihXa6ZBWJAzDl9xUEi2
ZWi0SYg0u9MePjYXmDH8L6mA2qidM2tjrW5xhbyk5yYVuTge84VbBgqDBB6eyR+8s2gM+hLBpGLy
k0zhgf7//RW9SzfivqySap226ljU9MGykYANqsNSAdf3N+2umHx+brJu4apgLNZQqrT2h2FPu8SS
3Mq35NtxUJ13h3URBpKNDPFhpR3Odozf/Ad/zT2h7Gpvn/WfI0IOjhqmTDBm0fTn2Ij3EGbfJeXU
ozoDMP1AStODZvUzIjpqpE+vcVoL9Ew4fuYLC1vJghEHiAdfa1raKvIMkaiytxQIH6HkmNzlj7sR
9PCl+KffaFjg75fYd6h1quCXNh5AknjFlEZK35Tnb7Mi7R/wWPFG8RdhZyZRQ3uVVx+fOg3yYJcl
SKJ+v82zSwQnzf0kggy+06i5lRQSVJKEcPq2yYzed3Ot/LVOwJA98H2oRdfULWye93HzNRPJwQqD
eU3VZGWQ3pMir/0Nks5GluSQ7Qx+OqDFdJ0FNkiNEs1K9owfgbX1Z32uapU1Zn0t7T7OXEldq282
ubwG2jrrkX3PlIaPpz7GhKFqQ4f8+t7Ytu5v2hCOU6fF/Ct9Yavg0wEjN0o3eyPtMwF0quRKAIII
Sj5bogRPOvtjHs1MckfNjfmbTwGFuDTIJM1HHqWUn/6Z21bupWgbLoOAMIUB4XxqlmAyHWH8lfqq
U6PzHZtn7vkoRsJ8sipqI+4yGcLa/RBlxZekmQor1XbyJcuxVjTYIH+3KE+3WquvPidcvs/7g/Nq
R8y2eYzO+39V3AsJBzJaqNLd2WCa0CytuFHQJ4fhL/nmTj10lH0rl2iyEQYlxv91lLuinbGHALK4
1nRBGFGztyEGVtWxzYayFUxdvHJFv7KmJog+F7ilda/ZzamaIPC+2lNLS8R1a1SRVPCSsIxKsvWI
qA2DxqAkkul7vzbWOwIKIKfaB1QLDEkAFSssNZiNEMnuxQv0BN7scdA38P0aTmZg0mYBut66bUKn
8ImMlHfkzJFvCA7Fk5lCgaxhc8EG/r9dBokN7ExCg8zaFsw6s9vFBzgXYG572hrceynLEIG0MHY/
zi3l4GttE9eOTI1RUWj+DYYagyNfRc17T/bTlD8eiyvIIl5yaspQNHrmPJcAO5ZB8JiPflG+x70P
0c+kkFA+JibbsP9uazhVwZPZ8x8PwTUzNVviUqc5N7ot4yDqiaQ7GxqYAgr4k7TswgaewPr2JuaF
lWcHf58KBX1USNSg10KboH8U8tsFtbA76nGIwPFTMqrH04sjIlwghd6R8d3AGjXCnV8omW3JSWMy
vZKtst6SPkx/hriDgV8JdNnYMdHbUBjFv6THISWiKbcgu+R9SzNwpX5FHebrKV1UFo917jBJSSN1
+UKrL3hKYsP066BG0ojvPis3tEMhGMOczTrnVXS7qbeCJeNmTq+F0iqhRhlbwgc9wClkEkQyiHkn
AKlDWbGHoTjyQY4xqoit9eIM6M7I3FI+FD9pMJrtOd4piB8YbI1BnwW0PDy+Y/DzIZQeaCxI0ZTU
SEczL9V8m8spDz6KM5Vsyaevuk32QiXfBItx8ph36iC3roFcfIsZSThy2KZfTStjtrAiEwRobGs/
plRyrT5yZQOESoVf45sjzduOlli4pi6LCW//OtBiAUlR+ntsvlLwkLql0odlTDmhhAtCxa+kxFgu
i8NvraRIS1x46FgBh691kOtl5HTIJzlNeiboGPIj2EvRCksf1iONdOHMEIdwg/M/zo9WBgSDY2Nn
A791OBqFYXmNzk9aGYYTPHTOgdLAABTBKIxnfj6hHxM/4QXFbApT/0uSJiS9R8kT7v2u3aZaXwnl
HHo3jl+a6Nu5DtIwv4hPrIeuA5hTcvT2r8R+dp4dNAOGivV5HmKB8/REntVxOJwoNbh5Xz1rJvw7
THtVWRa9dI+tnWCQEXEgLklv77Zh4HvKSB2NaHx9LgPAi09RxaJC5yME7HLuOuL5AHbWkj7V8+JY
m1aliBmP18/YjSDYENRaxKxbG1Q56Klci/b4dNSC4arWReuZzGrAfXDdrrB3NVeIHA+SnhBAOSSq
ehlz97nBduP42WWywA6iZVzr9SFG5R3SnGvKct47apchr6DIHevHuapiXibsThg92ak6ZqLf7F+E
53ge2tBGDLANbaT05zBFTWPvbJKvMKoPOQb0P2GyGksoJm63H59oiK+X8p4+aVgd03aa5vPmIXPj
V4H7fgzmudaL8KCfXlsVWw1gwHQEWUAR6dgLltO9jL1KZVpZDErdi0o4QHUeuVwBrST/YXKZMNbG
tpsHopvWMZ2DKP1sXy0++onQMx5cOP88PP3f0HD4/cYc7lDf6R42Up35DDe1KMIkBDgSqj/FUEu5
UWfinW7QWbx7seWEdfB2fJFe2wVwTGvIHQ8LgQRREp5ZQCwxJuc8jM0U8yAmQHxSyoCg78z1QM5j
XSGpExCYYFk71syJs26PSWBJKc+ZHuKQcXz2TyoI/fBacXZF8D6IJWzR3LIKjXvqZW7wIKBb0Qj7
i5UALrekgkM2ma5Rr/0u4ZdND3SToPcn8w2zK/8QWmndHsZ+vAKFi+0rKaBZc0uixPBdy3DJFcK3
GnM3L5Nes4bjkqd1S0PgSuksP+JEc01fr/UdkQKZ9ELkBF+u1PAEP0tcsXZTlq0EpQFEaPqHI8ww
sX9nJB0e/d1oTAkjKCtWlOGmf7E80+RRC+jYMGBZEJCVdUdSQfdJ1CW5c11zSPx6vIuLrU6oMtRP
YZBfLGp4a2yQcbG4Udw+jQCyg0uybCfS6pw8fElyKwnek/VBOGDXydtHXX+64RuFCH4QAfSF2E2J
/LXnWULOhc3jKx3Peczdbc2zPRHwa3EC68lg7Z+T7eAM/YKdmVSm3bYoBn4tL+NQZhsX8ScPHtHJ
7JE36dtUAXy/b5yyZpZ+RVligfeUhVCe7pIcIY7Ygu2W9y9c0f+Ch4EE8NKlmwXgDjva6WAiPimI
71YRkA47HvYrCZuo79aWlDK3oskWbxFU4CPtBFYPPj5KS9MQzmHkThpukIpwU3WkbG/U9JK8ps8G
Depm7DO41Ir2yKQUjHmubmN0pc9gUZmN58KVPusvJ21O7U0yDhDGIDRmtwEy+S8nrLxrmWgszROl
g8NzRpL/6o9L6jp0FzmPcX25xFz/6UvyHdhRHqyjO7CIJ0MiyutntKOSSrkvodFSjA+QFpbYn9gn
NfF8ZsEgxVZ9WxwX/FLab1q3zK9nMjOuxO7v33C7Go1H6e37Or9r12kA33Pps5XEWPVckPMjhERV
ck6zimk2BgEEhWf5B2LAomIXcFKQEVIR142TsrjV4TeIsgIhBze1rLGmsl9BFRsDG1pU2EdoTh9g
lM34svmDu93RGKQxO1/j1MRjyziX/suT4JHcRcD2eZfInTIaoINbeYWhe75fgh9nIT6xSPAEGgwl
WgiJplLVdDVg7rcHbGY+X+mlOVuMOXqO7wn5wIdkuGCQUy1GrvXUPchYoa0/2dPo5DbTh9mETNGR
1hSYuqUU71dbo3kddMpwKT/PV8s/NbmZ8AKqutrZb7YRwK7995TmZUztcUFFGD2qCWdfYsBvI5/2
kACCunJQ+YRiKsRQU0ve9uJkmPzFEIUSkgbpy9Nf6AtcQDbS4jClVloGy1wyraQp1ckjfTUz5zlS
yTfRZk7lAk4oWHiE5rIlxbcbHwMdJ6X3DrvyzA8rZJ36chQXH9KgO+KRPxxvO0K3IW4qvqAeyGOm
chO8AOROa6tqKv3xxGjlU0bmaQHgOouc1U0XpZXipungROYsSkjIcsWq+n7j6lsqd56Wy1+ygqTD
yOH58+ZY4njNlhiUda20q+2srEvLy1z2z82Q8loGx+wCMk+GNq7W+qm6X4gozB3wPxr+d9gwhWYJ
sg498alenXOdttbTiMrZ9S4o7Uu1vcA8B/cwe8D6KnizdJo8LMXQkUrwz2Jiwha7HMLr+WaXR6Ip
Dep7yvhww/yMgI2O1LPxueubeebEq/BMKDANaDiYs5PIuHo/bYU0SATUsdlNGFlH4iunADCQIFX/
3BKPQov3NsCpO1ekLEsROEnf+dkU91ZsOqyfUEKJjyDIMKeLrgTmsFNSqwJibkpU8gmHLozAtkwt
8wjqHrYMcSqWfOv/AEtc0bQa+ZLgDA2l3PWg2P7Igf5C574RGll+wj2/hd1b0Ys0f0nMnJspPIru
36lOArYW1Y+k1nLjLwag28j9iM+GaxV9oYtuNwwBsYprmiRcQuGi2fxuWG+Jyw4eZxrqDoUAg7zS
0B+dH2xBI/1tX2vwBLg20aQBQiwtUax7vGvP8BViS4OBUyc9njCGCouTajZZLiiCD8Mk4qh9VAox
HJPOzYO3iYeCN1A+lWJcERHSePSbzFpZuWyOBDasmhjRkKsmTvUHx33AihevmnO53xZb4PwyKWwU
VLuFdZuWfT3On5zqKbDG5IwrYpTRQH/3jMR5zi/4wBNEK/P/2asKibw4mX+hgnceQBlsfzFpEA3e
VjkvutxJxSR6bDmY9lgKOywHDjFzcFB++UewaXHg9RErCvh6y/ah1wl9HVr84GKtBB9DFdKkXDss
moR9xtXmWlg7tRxHjgf/8P2Qecr01BwebbdDFCUf8SLD1MtsYE/IrznmGjrW55v1AAnbhVpMR+cd
W0IVwYtXUi0EP0yAu5S+Bmr0KzyG9A33XJn3ktTT69jAIcWpdBa8jh2MDHopZ/uBkj/Apv7WxCSE
8R+lyP74LxXyL2j8MgQaipEip+ijKwHdu3ZDrt1/TyZukJBDORPixOMF3/foNyoIIS30lIFu2TsB
8ECw9MUOkTt76vYnMT177Yug+kXA9+K+z/caYFKDbOWnbyrRq9YpX7rRZfBU7b0/q60si47eKlqW
cGf8znrnvbnFB1+YAb6omLQbd8n2nprNW9UiSXCrJsGFfkQnsvysNDBlTT0AVgLZEIbWvH6UiDNY
zlIdiArN8mNrwA9ffZ3SiOuKTiuiSnMNvCggHSSkMJPsAhEXNWBaAsY9KwebMUUmTgNxrW6sa6ug
8+U6qrMVZiny89i0B4yWS4hS/wMfUQRbWRYZk2K91vBDXuJHTFnDBR88kE5CwVDjxgwksskb/uPE
JXhPHgGtEvwfhF/xw2BqCbHDFXj7YGb4TC6UNua60UNuyI7wT5TkIgWGqVFJWAJyB1/fg8CQ6NVQ
cB4QzCyFN0AAfQfIb7vGEi8nDrmUbooOXmArUJYeTPjDGl46KtPMdmJHXiZnLEyie3FyMNbLe/95
FyLjFrB5PCzpI9Es0XlrTseC2a+atHQcow01amcMhBl01+3gHpW5A8IfskEjozOfxulYpwhWl2HD
jYa0bLOq9YBcKTTC0uhmAz83QeZcGNY5t10+ICksitpL/JxTymnWz7ybuI/1O+18Rn61EK2eXrjX
d3E0Hq0N4MIfrBhQIOSzlmSarU7CTp5gDpqUKfRQYAMeiCp7Qrq1cAprPGUzKoJbBON9eREtAPEN
DR+K3Ok1zsO88o/ScEcKGbx7tsPNPWLSqyj5YyuuA2G6lI16iK3PprGFVqohxm6D6Sox0PSJvC10
TTm/k+404k5AEelTuNW88EMlT1bROtlLy5MC8nVysJuPvgm0P/huRHbc3qsEhYkKMbcOFBD4PF//
7Yqbb1W2NGuU5MN2lfSV2mxELFhWqik3AjDbUkxfsGGjdp1fBoeq3IwpGmRqiTgOG1+ywPWglERg
EthbDR8I5cEaAybeMAVPzpcyvRwc0eEOMta8A+7+E5BJZq2FCb4okneHvQLle5ydnU1BfaKm7aCN
FA6WQj+SoMMhJ5DOkC2CDDNJzNJuIK8sAQLUB5KgGayYHCn1zTVXWFeMmO+U2wsLAuksR5KSTtST
4gfIZxBASVWnnJummjEUAnU62l5uotUJGXFTegn1J9L+bVPQgDfKfgNDoG/2BkbBPR28l4QwmJve
5oWzV46YRhSDsQ1J3qwWbuefw5iBg1Mfb/3h9Go/RrRVTRDQYxPDqXvPvl+P1eL8o7wbjJ6bSwiN
1z45p+LQJ2tD+WzU3jaJc3mT+u9LjyU+LWdiroqBtIakuVvSiKukuv20RdYWEgo15zmZVgQM5lJ5
PeVevnzUjofNUyJTEFvYi0eCBXFCGOhfzbUoYMLuKs2WWBBoElZhvDdysWpdGJBV29CeInWEApqW
Y9sB487LXudN2o6gjCLEevBepNEM04JI6Q+efR4GBNVn0PgEJuwShK6cybkc0ACmf50046duyJq4
kFbALvmgjDx0oBKAgJWKjkdq5WMFm+ck3CZmfgNHUW3fCB/vWOE4Cd9zau0endv6SzAxDHKWYxN8
ke+bUvhdpZXqVZeiUOSngL/ZximtOYubbHEBqii+i4CuGOe5KDcwm4LVq5C/qM7QA4amnBgk6wW1
zcqb0JUmhxgWXdRDbWn7UN/vmPMf5dVInfRrZIIs6o0XAiVMe44GqFF10dDCwCe6g+TxTIutPqHN
xGTa/cJsliWRb4FZDvWrt2l6AHCAvV5Y54wN3dBf3GetHQqdA9tlEBaI+MREguqoz5fTUAoGExo+
Q9PQsW4CWTKbMUMfaj4BVX/uramer/G6X6O00UqZqCLtPHJvM4DpchyPdyTCNQitj5XA6A95xAPu
laYID0RS4LB+2R/RZn3ve2gcnUUV7MptaNyvJLDBviNGq+X9Mvw0BEQSNNEAcijVfErJ9IXtc6EX
QmSEA8yRcb6BQfe0Xd7U1DVtJG4Q1FG/jHuV6hAOIGbD6QEGFUHYH5ZlCwryG0ICkVgJbFNUGJbX
/gBvZyMLbqFCYJJ6BIUbdEqlNlWF/TSl0L9M5fGAno5DTA2ZyoVjRNqZJEkaZVoHfxynPQZbWvlf
JHicAy/BXuRRDv4ykM/b6Iu9lmZcwSFFFvzng0m73gajrcKTJ9yVJHYk7TTZh4axE6LqAij174oV
kQMCGUCgPsLQQGC1tJRc+77HkGaLRRiCbu6HUSHWEofNmI6x4uoFsA47m8NEWUlxRzCwWTHxZV3n
191GvgPFutTwG+dVMng6ktKdCxEU/YAfhkHkDd1wA8w1AWH5lElFNnXKytCQ9T0IzWD298b6kxaS
qY7MuUcV3Fdt2pGqEcPlgc791jonqe/lnbFKDgnoRwh3hLUMop6mHkr5tQS+e+AoqKlc63x4Z71/
N+Cs1MaxiXTqIEGcjkrQBRD11JA0oKS1PU2MppbFIpzTfltSzrBpPSwfC7HT8kdQaJOcEUr+YVrp
NIXB29LCbr81S0Bl+BCTHoM2vA0+AdJFS4zh+iIbEK2w+76b4JWspltsA6Fk0EoltqB+fWdngW4t
2cwHkTIecXQgDBE+njX85imOqNFq7QwCt41kmi1pNSNOtX5aLHCUUY7G56aYSnfDPhEvTOrE9G33
87bx8tFpqc0nXpgGJS1ketgDjbFAtXdHxYvjCfQnVdQ3jjB/dcGTcZnIjcFAaKYRFdhG1s4s6q4h
m9K+fduoOyL+a1uYtpjc+TSgs0JdE+vUjqGoAWzCfmLEUagfTzbxNMc5xnaZjFCG2zkcBSJs94Ic
HSVPnvielnT+Xp06eSuRF767pKqC3jFPG8oIY4LfcC8tLLeV/li4Fxq2KTm56s94duXRvvri+kfe
YwAq5+mkj0rl5IPUbkWvJSTVXF+aTyHcjah3dvUbxkwp1+syEoIONxgCZvoaeO3Qwj4+5g8SORnq
Pl/xYScUFSGaV6GwyIiua9FMyDlw4uc5PDN4Xb2og6v1HbnqcD1Uhd5SxDwySgqYrBC4gHgnGlWp
ZuJrVm4wW2ObfSFROm9ZCV46GeonzT9FD495CMWXtzXM2wv95AbLUqjiNFJkYbUmSeVF1/jp719W
O7Bo2+5Hs2vMjZL+TbR7mCjbBXFfATKiYvyaJQSRbNN/AbEa5NbZjs4G3sxX5PPYVSvMywO2t3Cx
weymKlmyfU9lft8mxSMR3J9jI9WmhurMg6DndyeUWorDHoDK4abkuFhhwKnWTn7HKsG2Us0PLBQ8
RUhcj2Fw3GMacAdbbaSW0l2zBtnax2Qi6xoJHUUgclSKC62PtsBxbpGUSpkNwqE3nNIjgww+g8sb
RCjB/wZ111NG69E5e4oW2h/xuKcoxteIFgNNsS0iG6lDsWgP9kgzOHke8sSXQBqF59JbAk4+OFXm
vzil9llmT2WbEEPXoA5edKhs/rZk10MKXatg++WjL0CVlJiKpZyK8rVfn/dU9QrR+1F7xMnTRTPB
glYfTu5ZDMbXcGPsce39EDXqLRt9ShaaZrD/4zeJfof+gRVTvnx3uuxkbZ07iROSybtFHhr/C1Cx
pwoJPS1aFGJXz08bClHRGE0Y/BPKNpDmE0fLnriIdeS9L+fcpppOXZCTgNkiiKgDzZoWqsXO1Ezh
skt/2DEuoKjIjqCv1x+RS8n2gjaqOuT5pcfMrUuqoVb7zx6jD17KwmObIpgW2UfNyOVvGUvK0jX7
rMaJ5v8MzSuMs+D6v7hW0hie8R7tbHlur9Voo8eCKe8Zy7Rwpoa5J2H+P5VPYAOCqPnqeYcp4O7/
ESKRbgb4AiBmHJnm48G7eUZ5tQvW4N3el52EA/gFBnkYvVd0jo+VePgGEI8jWUC6jIGl1+CapjGH
ymDENC1FoEBRUYqatYeLCEVdjkjX8KN/IrMuFUjym+8LHbcMcmsfK7TvIFFoHCvwJGPjvfPV1l08
NOg4DqvmVOceZYGZmTThrBCOIj9xfzbwL+HEkhjotBUiR0i/T5RKRACo1F/Qy3LGKwigEiy+ZLQd
AbfHzbP/sMcyOoQPeTasHwVPSjGncWQHi+KE2o4Oj5RsmKK/Bp1X80abNqZvTqzRQOa+5h0dhl50
P7GNhoQIiZWAy5WoHYWxXzjVCLH7e2F8ff4hHdKsqmeGSWzdLlHdbfcrvRSG8ZGPbHBsP857OSeu
ElcsOs/TzlF4CCuRthVfMWLpOTQnbq5DCsh+CWrlQqpvfIJ7NtbNIyuE+WckKrcCSwVlymRfxhV/
f344jd3y+nh3aPQSr3+FgE2agv+9XbOT22l16AzvVPMiM3HMN0k2WJR6YicLiKDhkaMIasvWgYND
BgBglClry6t+L/bNn3JIXb9LEiBPx248PWgbCE55R3+YxXOK95IYx1RJ2StizlyyvjsWcOq+bw/T
rrE5c0WvYPY00MGk3rkOL6k0kqsrf9+8B1lq3aJvzi39wmzCODSuKOMC80FWFSc3howqTWJia/6F
NUpbdU9sIdX6ltZDHF5Mzg3/rvNU+mIcksRvCVst0yZZ5UYaXmFiQOtDhQ1ceEjiZFBjePiZ2kv/
ugOUs7DAV+ROtjQw0tWcj5t37pQS8lP7eFDiFJz9+6wqLnyvAsqeT0uPhMB1di6Sa+Huhq8pcz2R
hGcx21OagnwlSay8zsH1ySKq5Xc9ZLJyIigpu056AOo0exkXRBfBkvD8nBN5B6ZrnyWEoVJKIaLS
Zv73NkJKV7SfgALnBaHO9wC6QxMEsEAR3xhM95FznrMVbhHZOBKdPjVL3NeaYkyrScFEh69pndDc
yMgIwdlgIkcZxNxR/G/KwMyJ2LADlxNW6V36z1HTvj62hzqMRN9orB/aM2mq6jksS787tI73SpJ6
daaZiUFbTWdmysmPtlBBr/hSlF1wQs8tvZz9DFOyUAU5XoZSu394jAtJlLVGJfwNVP+VGquQAgIT
7865xfWvp4IFS417MkVHVP+/JtuEwPRMRwo4UYLSR+6XTJh8OZxTtQH+ilEFzREret7xbJYf9N4d
HJ87ZhkefxSQX6Za20A748yVqnB+gMDX3iCi2WE4nL5oTmEh+HrHoPnCKlQgWPkqFaJtOj9aPXI5
u8Geluib0OA/JCvQnwvyuYqWvZ+0XnTy6zkfMOpxYUag4c7q+fyJW2HlpDOCrKZbviIZASSkrTaE
60LLJUC7S398HJm9ZzXxYjJRglxnHxOpMraWZxiHmtAEDR5d6eBblKaL66inl6rjyL7fP+cAOrDz
VIK6zCCyfxAr8Twuw2rr33sNXBl6msY5G6c14Ddq7bZkvvLuZtJg0nr7fqhe1Gwh1CSG8oSMf/VQ
sGgdEMriop7GjOq7OoQ9QFWF5OXB4EAuMc6cVrA7ixFLrePV3RD8mDVL2/DKNdC2ReZ37Hd6MZJ3
BSczqEZBUDXSJHj3/T33RK2DVo1WJMFgvHHcAg/+ZkWq0X0RXbAb5jC5VSem1ibEPv/snVRHQrrr
qopKAvrMA5DO6nd71lbS8gyst0EFD9rAkxnwUHI75rRlHE1B7uBhAetCpKaftHHBzqvPZVvQ4HPt
8xRZLdn4QGfTNcfOpKt4A+DEblJPl1B1zJ2vt80+fNPW4BB66qOWarGFGTygT2+kvr7rJ6CKWse/
dz38cis5x1AEzpad0LV3wom+4Y8YNff7BwGEq2CK95Fzz++EcpqBcS92TECzCZnnIc1y38ZkD4rM
p+P4MMd8I9KJrU00DYVOFfJGlPugmWVzPEUjgsaI2THEercNZGHJgPVOxMPJ90p2Nnk4Y5RPqobe
Y5zf3krmebulkAqE/+Wd1ZgA8xVp3qpOxhNum5B6d+M3eTt7sytyJs7sRTi97mr2A9wICIreGvO3
SRaHex00g3HJMLZoSeWxz9jdxYjkoPe61+TL2ONRPMYjRQviq7hYyuq6gpXLCVoaSBAb3EJ/nib9
YnKswibNvrcvO4vDn+s/8qjDyW17s5BN7P0yt8gcRraQI46tP31hNexarT+mQGwGP8Vywu7f4qml
LfKjD4pmV8mtFIkS8BUvY1xlzfVgFSNkvJPZQhMvOWbSaX/GojjCeeFEvpEE/xHKNduhwtW29Adh
yghH1RYxSx9JTY1eIjqfxK+ynp2vRuDV6P6DTt35kEoYdNc5OaDROp8If+k6UEoAuAFgP3GmB2hS
YlI1J/2sHQDKobZHOiJzkx1+MHDFE+FiYTut+4vSAqhO4zjv71YYdIAhQ+PpMR5JdutXb75kgP+a
5VqSkruWP7YousPNFqbd41J/Tb3VLbfB7dDtHkkK+n4W4+CxRfjBLWS/p1qPI3b9Cg97XLwEfo9V
+P6JfkpJYq2G0mVDR1PNVR/N26WY5ixd92Mspl1QVdM3bZgaKa5OiKk8Mun5mKGUEdGB1aUvW/qS
UUGU6EabOIC6xpKSI39e7sI/W5cudjNReyKlWzRXM5YiiFIdzPJQg3lNrmqf62YyTUGu3xTZw0Xd
o0RjATB9ZDjGi4SkPpFIci73q+EFjzYBB+esD7lgBWhXssMDSibFkF+yug7fc3pYB+FDwa+k+ekP
HoWysufiEHYmmY56YtKenD4CA1c8zFiJWjasWjbCR+UKjfDqsICkjbbbfQDpD/mt8B+eOTMTcXtY
cIJ0yL1nvE4nY2wPuhNw0UrdMnrYd0c8uRoECstZqXJZKoVN3sjrQkA1YwQiSllFv4JQbZ5htGVj
iZOKgkLJlYqTHzc2FVU3prl/byqq8Rm+wY7/FezPXRfXHNNq29h2GNr66Ya6sE3cGdt3sQnKMzsE
H+H+HJfJ33Gf6pqGUcgs7XCNwKqL3KQXyZ+hzFTHMaG6FGDFdhBzoDpX7mJaATetnfKU/TvvL2P2
BRZo+PpFlfU//lO4i0nMt0uwFwDLo8EM+3HANT9N3uBfPEC/9e5ucsjPKYYOQgqZfpBx6xR0Z7o0
NBVNLK06Qn3Dxfvek9f+EzY6ASOvqTdWK/FI7T5ICesTfJsv04jPiSlWSVei39Mt4IwXUpvLl2LM
n8EdzG4md1YEKl5LL5pX9OiR/HN7nYfwsKq3b3XGiC3ESGanuDm4d7hZu9vxe9UJosG3UxjHddog
HvN9jtD+RmkKGSh5D0nhncp5g/HtGiAibUQVCid5BRgj7CrTX2Yr0zgV6xaSlhyZte52cX8PHCl5
EAFOOTH0PvZtF8EdLs5wdemH3OYTlrrlpaE1AmDRhC7aILcSmidOY+JrQ0sk5eo9RGmSS1Wy8mcS
VJNWv+O67ru9y6OYxMI62nswluCVvwYrSvq3B603c7PxX6MYb+R4on3tlX9zZcOOQOBYasYlMkMM
PGvjI+ZfpuQWtb+9leKRXH4VgNvIX5HUWhJ7QY5AiAy46+P0svjBhsLkPD1Iev/DxHF2LZvJXAfe
w1GbB8VBqR8hi7jhN0AWJXZvyrIn3xnjKnFMYPlutNO9PDpd3TgoTwDXXzd4/VpS7KTm86bfpvQm
BA82ypFUwpOwNhWyoHy1wTXbeysAdCQC7Jb3zHLUkQDX/rSD2490w/FCdAns7+jHTj6HDqfntJyd
jCJDaRzAbBTAciv8gRDtIcMVWFhH3kQw67cTORnCxWwOmVWOAxtAaKe3cgzFvjP8Vuhtg3RQyU94
Bz1EfWHecODZAEezAcOgrEZvAealxfUmlwt02khc2zxR4HD3tDfQh/ZWbufoKyo3kXiLULYE/uRr
ywfqImB7ee6+h5+u/1rNfKXWZy0nUavsMsuyaq8kJZbzEX5nJwdso4p6gP7Tq+/uEGigg55jvFh3
d6MKRwppID1i959Sean+KZV6ADsq/Us2HShpiWAGmjHqXavVRH1Ku7wus83vSKRSqZYAFDNu6CYW
sIO8ZBXCWEjNKtwa/yQKsnpZl7GKQ7ArRpx1QI0bI9wPQ7I49eL3Cl7ha2TwPTsMSKz3Tab+6oaI
se9VMQLRkGUfU/K2Zrxsp4S13ozlcFXR7hraunY4Kobx9C/hjCtPhcRHtOsCe6IiLTOkdbawiCmd
h3XwC77Dfw19mtCo9RZKtBbNj3tqHXbqmkK4xVSua8SVnCJE0wEamel1GqyzQ787e2Huhfz3W2PU
ilNqrIvraq48xwAvJGg4TQcC2f6VULSqtXr873p0/EWVJV6lwcFm98iYGxpDMPk97rVPzAL3ZzYS
nBMqtFxIO9JP3LBumtBuSDdkoGwyknnsAAHncqtYgi9gzIA/FOwdLmMoQQp1rsW2hXQwEA0v2ROo
bZfeeY0I/FA3acIuAAkmfUD5ecpAow098DrVRTNKJA04dR4YyarBDJ04wjtXoeUa6U9dT3FfIk/p
egZHtuan0s1jFFxNH1UAIlaVJ2THbJM5cysSk5UsXaUftH2SxGGnKluKePBDF7zt+Msklr7aaVOA
wABKOsx9DfnaIKemmd9QjT/uWFlZdficQml/zwNNi1B7M67zlOjs5teGkr+6xYp2TnlSlMGe2QjK
W2VDHTnhQviCouze4tNwqgKxP+wFNjHe3yZgzw8gXH9QB/kPNBOjpFotuchK2CMcpxMyC7pWZDbm
jAdPARjdiByjfk7TgX8uHB/Kg8K4nwu4VmKOzM18vxV+jqza9izXEbN8irhe9bQofUqa8PWOUl/3
5PRPXDRQ0s62Eq9l9ckzfr1V9FF8kF8ViXR9FDgfAnMKFz265zADrdfDqM2r0d/PCjVNZz0EiDgP
y0+oNGkyUuOkZmcwJKnOGQvWiPA3ZVwa08F4OSP+07Pbb4kpf1/g42rzDajjbIyRqNeW0af5FNHn
dRcEJ9KgKMuR59APFlhjUKmgt5Pm7q/xtYZwc28JtcWdWO52XvumdtNq7BIdJVqJXvSLYVzBQenB
im+WtoywLSQD8NlY1z6IoVQYOoeooxJ0rlO5PoVYFZ6mYvKvd3BYyOxNpa75ITMXgUkdD4rduWlQ
G6muw2TbfLowxcF20H/np0/AmT7bLqoAePjelWwt7aZS+X64v2H4DGToNMckG4ky93FXtLJGiuNj
FH5N/KVoBrC9Lu9NdiQphyn30BrU9HOz0I/QH+vJjBPtIeW/iPiiMnJwNR5Y2Q0GSt/fWY6qTx0O
y5yJZJfl9JHv/acFG+/AOWCvxgQ8SGRZS7LFxfgloFMW5WXB6RR3FadF+1SgbJVMWh1RZi5VD1Gf
N2ELx0GuGsqP/7A0soleT6++agyxRcp98ugwH0YkDnylq1C+wjxk8OXzrv3aWik07Hyn+OP4YwcJ
Dwmtk/Nvmw/FIpSgMwvPUXcpPjy55ozFceGG1rczRTugCD+4IBMPHJVzlvxG9B+QZcqwuDsFwnt1
r4/1yapzN8OypbtBZXqc4QPfXyt9uLCI/CjXSnAcBZu72267R8+HJFgd5M6ddzzFRf14uGZckRMz
1zJdjVlC4cm8y0xAJPIrmxfhzWO0mYNnBi0VOrOr/zMvausREUidwUmd0DkIfjAVKdqiqF2wfbzw
K8wWS0odpK0boWyZ6KHuejdda3c9a1BUClqkRP78keD+JPA67dKe2P4A3d8yVF1ASdjAxP3q2JVj
43swtsuO3+QekVWJUm9mm/gxCpeUc9/imWq2eA3OV1Bw39eH7k3jSol8IEzqhDVOhCI/mDmA02RO
ZkA4MgKCz3NeOOHr4i5jgzVH2kLjL3oU+raggdY2+Byq+0mkyctxeKWm98RubawNkMZf17BqHDf1
pLO4uMrS62DXHYoWmndXKCv63/dnnyUlq+T7qlz9RpRFXd6RqJRcM95LVx2v1A3tiyK8RnWbXa06
n8smL6c/JiMBCcOLUUVysHNv3r1qIxzrFTUOM9evXM8S9q9LK0UA6Okq/ALivr5wwlmlhWke7eF7
uzNJTfLF4yi4/H+1NI0NVDyGgKNzo0QUEeEi1XXj7lpQEbyF0a8i/St8lMidTCl32770F+omGaLF
PssYiR+PDXNh98n/0fblm1e6F8L8rKGun2tuHmgu198lRa+r9+PGj4XgAZNBjlwmxFObivuDpVhT
1/fbeJWBTudsuFZWNTOvRPt93jj/vedpRhpx/feyjkrRHlilrtjZWLso8Ck/7PDf44GTTr2X/dVf
DLwqMqNM6DJTD6UiKc3i6QBqNJju67ORi2LM/SHfZDAuO+LO0tD5OdjZ/f2eujaRL9SLgpnzSYD8
hvLsfM/4MqtGTWFj7NRacx0dRpZgFsgZOavSS7Umtc81XB9WwEfhsjYRC05+DnbZqEs+bA3/D5pk
miUlGk1UWIL5GEL+Ml8BLSuXcpVNEVNGJE/0Bfh34WRNCP93I3OpfB+3f/YCrkAVgRJ1WlthENRd
fqtmtAyVnOza8ldv9epGWaA4+XZp4J4DChMd/M8znSLQtUniKKxHUriZgvG96yKmfycqjRUJJ5sI
31IDHgSTAGO7u1vayolp0Ibx6sISIA9xq1xH040+aqG55LGJw9wO9LnuAtT1E728ci11xPOahs9L
W5Hj+/fcW0AA/gLnbC661e/IoksccsTBnCriwVtstNJj8UstKQQJEgk3XhuXWMAcjL+6HB3Pa83P
r5JxSJ/jtqGKaeCZ20kGCJia+4JBoDvgApIms2dF6ip8NYbxRR89NPuga7rRec7+weMwq+TUiSGA
LM7El66F8xb80DqZPowPGhjflHBhWz3/PpkmkUwGuGFV//Dx3W7eX+OYMsKD2QNbTwQ3iIeJ6fl9
VAdy4Gv+rDXDA3q090+D9ORoEtlQA3WxONtkT29hILboyMfJmdiFVqjeVHxb2EELR7bt8LD29QIn
8rE9uVCTQ3ReUsYD9SaFC2hwOsOtRMxZbXTaRFXGPlMddtvbbrNizXVH7wwHmr87GL5cpaRzICg0
AlJHGqLj9ncvgsxjny+QVewHvUeaKcdCfSPfjceN4sLqDCsMKAUqP/TxsMjF6FJZ0Fiqx/1XhsbG
H2OcOR2C7NMF5rSlG+oqIeyawsgQRuN8e0T6CeQzxsXQx9oMDsIiv7m1aVqlhwzMhh42lXMrxcKH
Jr5UMZXsTyDNscB1OF9iCwgWDZLmsS6rfQSwNpWYSpYsOP3YHB+6qokHbe1l6noOX0zN1csrl9Jt
I9eySzNhtyaEsFGRa4sVjn3DHg348LfIxkxOkFNzVZ0gVFVX4mmi+oXxXCFMNiDaoJbZVEq+VPrI
tbLvW+pXWMtbFGV6c28XWUg6RgitVnZDbGBQxBBqsr68lrrkvppAnyF0z/Hm7qMZe/VqbWueIRZQ
26W/GYgDr753NWvqn0ywMFmEYTU7cBAYV6Pi31YeHl/xRPkr+IvouT4vafdc6nZaUDLthjc8SGVZ
/+uYcYifyPUxZWfD102Kff/2M6Ho01hvCWXK/879hTtWxz0eXs1Lw7wMngrgUIgU+QcLvVEbB6YS
KN4nH4I8emtC9FwmS9QJVbIRlXZG2VEREPG1BihrGiSE1qwuH6vhSShmDlhnJz3P+1g3F+/vzSnD
/7lTBqLKsSGWCz8J1L8Ru+b1MKdZDegPRTSALS78tF/M8vS3Mf0PeibN5fF/rN+YSFkomFRdtU37
tpfcQe7kj4TbMBYBEymgDXYtybqKkWxRW9CEOchKK0XYx/GWwRqzEms+kAlf6FtijDRxJCRMHmUt
AvmqJj6Z4Iv1153h1KK7UEWCNt5ohdHkvixP9Jgzld7arGp5u+KnjPriHdpweVoW7SLJJbkS+5KP
JL5l2y3CjKgO4NEqsiUdwi6z7fVtu0V3RaN6D1/tKgxj0MJiCyXYincd/pmlNIt5Zw/iljHSTLPJ
yes2SCQW/Na2bNaIQHMZyVl8ayH4jiHEgpoWaiJ1QymnszvksWXD1DgRRvs6OdoE+MBT4aW2CNIN
CQYaFeWXMRtkxl3CNYlM96ME6GseH95X1YyoHMKeIcTRdd/S6WEVsCMuO2LYT/1TRAJBlPLpmchu
7YTLGaYdYE3MFcMwbO75KEGhoIOnT78mBOJC/pmbmNSamX8ZkHTLeA1l5E2OBp/dEF/UbNff8bc7
ymWumARLsTSl5qqGdT29MXgqnmetL/AtJ4MV0Zr5hw4CMgUMBwHQRSYAvFg6BTbRF/Rn0qPpn2Et
Y0I7zs0ApHvRgqZLxPIpVJi0V+CiHWvaorJ8husFw0CoRmO85Gu62irYLHvg7nW7F/8dOXy+9o45
TXoNoplKer0iUXslw9LSo3pQFN6XLxh4fV+QEKm2vE/DpXZhK3k/TgkkGP1609WYx0DYAY1raHL8
Ive//X956ppZU0BAMmE54/bO+g8aHqJivwan+cqrvpbKVZp6yk20P2UVxXRstFbrPy46Cdm7OwmY
sbQ78PrCOhDX7jcVhRzF2pdbk05uoR6gL74AdXqvKwI3mHcVA31SnjwxhJCG+BfMzdI5WOtelIMa
C1pIarJvwglcETuQFGjyMVYj681M1KO1TUQCG5kf3N6Xg0VYiNcROhNmN9LrGZbZFADijqc8yrGb
o//zhr10l2JUjjMKDS0zH4JyU9l/AKV93AaJsiVZOQ2IptEmazdt//kkRusc42xnGPN4eUDr74F1
9zZtiP3Hr6q2yjFxMQvZFnqVdy4LJXFRsIdPvoocDVY4R5mGa3jhc9kFuCIBRCgQqDHQqBAzB6Ng
vhYnZncUK/q9q8p3rY83IYDHVnarQACjJ5ZxiqUD9wQU7yj+O5+Z0SQ5XogE3d549zh7b4FbKEKi
hDNbn1NaFxBlb+oBXK/cFsE3fgPeHSfRIPkv2c8amtERjxM4IA8dJLaX0dcG82/QAZlUpyOrgYx5
feC94nbrZJs5Z5DV0ceGpxaDzKN7hYliyxP6hWsRgvlNlBj0E/G7+w0j/x+FDJEOGpDwayHbhNUA
xfMmsjx3MmQpEU0uTYyk7oqoDEpZkztK/gbjNsfhHlKSsI1Rher0zxTbrvBjI5FbQGr4sGfRby8p
DRN+cobaHz6QSdnSCnFWy5ftXHIAq6yNCGh4S8I7wKGF6msnX304NY37ylhDjuoQiCn/BYOToqsv
gcJf/pAUt06igGSC2VdvTRQjMYtcAWBVfeiWNXkgRPmU7Vi9lcmyzuoqTz0Ja8jmOtjUg2o6ud3P
q8gau5AQBI4uJWmLHAZMjY6Yrh+QIpXCTaSDsYMNmzP8zEHf1mSZJ+V3MrhEqFAI3yu2SeBDr43l
UgqJUW8bAJwn+hkR1w4+GVAehwceZGpHSSh908dw2f9HGoztBYszdCAMuiEGv94LPqFrBAM3CJD0
ydMKW5yEuse5uP+yz7Yk69qWoJOkIxqpsMMwt+JqPTBI/MAQTHJTsIKAuIPZFf9LBWk7fqWRAty0
tZLxVZECMQns/OxXfGLcnXrTK3eM9SUpcDKR+VmzQ+AA5OV2sPMy79jVthxu0Bxb1neRn1LUTb+b
5JPIRaPM8q9rFqkx2KaD1XMFPTYoWrtGlEi6ujJL8h5xpGbL3MZwQPeUEM9M1F2bW8l8TRHo41f9
gJTYL8QxJaDHpovmMMeqqug/C0PENaeo11tFCERwKbxqYychw+4LVDIXfPrw/85XYeZqdj3Qux2R
OsBcphhxDJthkGFwcYaAhPrWYae/5wMqkX6jZef7hd6BPVzOyDPHsW7dXL1HnipPNLCyifes+cv/
mY7R20tIq4wLT8WA0MJvFqH3Y7gy1tyX4qQKaUMlEQqyYbb8TdAWG4la40o4XtED9KL6tYFUVL+3
Un41KxzqzjZWnPcxJda7xp3DAiaLHtTzOqk/torkijeH58DIijBtdyfldSfebz+HhUna8hvxj0ld
0FjD6CIoA/4BM7/pN8Aadqk8TUYl/slNJUaZpyjhd3NQlEMs+Nsau6hF4LCOVuxnXpPd20hNsuSE
77/GIdeWcmJLrRGtS1h87MZGZH9afANbrYZEv94T5S2RTwyeI1Y7cVkuqjfBGn/m1h1L6yPqKaa4
tvvdi2NgqaP+zctKlIaBVpzPTQubWbZrd79nuY9vXB/QOIVXFXjFvFAFpI9bTz+RQBO6noU2743t
NrMuEXB2w5UTIOwL/2jfwHLB0KBuixRtKdwWv9qAF1Bu9TgZZlCkZLiEx71yn6mWWYeblnCVUDrS
IzMzdx/zknYCTAJrjjcDZzcwpLeU/Qcu75ySXbP7uw69e+Sazr/glYS34nSWrA9oUNChUhky1Hj0
VPjrfDAp/GKbf4P6NhXrWqbWKY2WxtX3ghj+cZTG+uS4fCwL6hxqhoGr/2xNuk9JAq2e/TAWCKUK
3Qo7mpQPa05WuG3VLGxuqNhpWoA5ORGMe0xLZj18amz5aTVIbfOp1Uy2GLpR5Ygc+gvIIJdUl22s
CNZOvM8n7FvEc1vKH00Aj7mZzoYbyjuYVk76EK8/LCEQasJY8OPxJrcBYJTHQ9LfDFZsgdt88WrP
SkXHQnOHw0ZrzNCdKLGkuDeasQ7nvcMv7y1KlekvbuGPsUUpTOd1AG29GMDEPuJB3wjfu6TrhvNV
uCIJsXmKztQJtDfOFyWPS+JmdFb4cBMoj9LtPIkUgU7Y9oYJ/0G7vDRdTuHUKS839twuntryD1AE
L7VpA3xSsBJu4WPQGMtt2uRwKf5Eq6ymUDTeOS5KFxc+VfP8zvMj/OKrid5sDsRzJLWcBS5EEqLG
pVqYYXJ3+XmlD5bt/YlAtCFEd7mPVDV5+eElNDqvKPmaM7XODcn2fkiZEdXknv/9btTpUmM/p49e
79F68EtthTiOqdq3WWs1I5sX9UJery8LemTFo/CUJM9idoXmTjNFPaGURBPzioc1VSIOWT5h2sZR
c1NzZTtefW/8mPNYUVdanA/mVdNfAEbePRqiKg/PBWZgQN3HQt4m2eopxH4VpsADF1TPSV2VHpOL
3p3qTk9HT+aA1I1BQYkcIF4mVgWYymnIuKFqUvK5kGJTRQyQZb5i1r4ekNY2aHADBzqvtgurO7N8
qSHrkF4IDHbds5EbZNW0ybQP/mXH5ur7Tq0g/yhyZ2bjmUEljFeQf2ufg8f87bFM7paglWlTlkqr
aTKTe972l7OeYBaUOlBpwFQQ0tauZ/JVpNAwl8gzRmoyociZHUFsnCHQdLca+Z5lYJ5NUgJ8mMTr
LEt8yCwo8GzwTh00tRDn+CK/e9aFSc/wdqN8lMbdyTGdZyiCK3pzX0veoUEaHTI/AEMQ5M7kemFP
pmjeqS/88y8/iAm3CYPzygVYjHtcvzAiKbvYhC6538bYdo6dL8wWrqCJdrrgSCPrXwpo15TcpSIS
u+4n5HKNgzcBLCFpYqW4YVgydnbHRkyITkdK5hJLt5uMttfrWQ9euqO9a9Xr6yAsfVw9sttGKdUp
b9K5EUyguKNh43wVav3cWGoQ30M1BOI/gry/D4CYe212xfvJMN+aOQuIh6sPPuXlTEZnEHG3Aj+x
lfbfCsSBjFutt4Cv0qTEGumbpkutQaARB5ROnh+AflDZLZyzgupxpkprNnelQlQCf4/skmGiCyHq
pKNoPHA2b2GU8dQmyXsK9GFmg5JMiv4YcLmg1DqGO1SnYu4S8ArnctKQHwfFw4IHLvWHeL6xjEqc
sGDL7gpoc0PiRTyvpEitBuu5c49t6cjjndtGl1iEfCKg4lpGYwy772+2dgxTVT+EnOA6KQrVXK7D
oGRtJGq9/Os6zf2xVnzG1c6SugQ6iyHnFQuu5d+TsnAY4+wRN7zaSRpyTPWrIx+XCnf3lfWMx8Rh
kZje4m9Q6cdidye8AWtZzP3YKI07FQOwT52Yzl8q+xu34e3QL/mB+7JNW7TnlMirXerZeejDHXNy
H4cs7hRcccAlmk2tIJdTw9VIi3A7bWMOi0Ysi4JM5gqke/bu/8u9My7vwPbPfn2wCYw7DdlzCEoy
X5r9DSdPoNp7TMdVT8TabN26P/aa3aFGx+00gA+0oGw+kQukXW8fnEPCaf8DIp1Q4j/zb1aJwK35
hzFCBXFMzb2m1E/Dnsy7evAV4h6MPiFvawGLX4zZjON5OTT2Nx+O8m6u/A2NtbgA8G35Brhv7UAZ
eEjWMH156axKn2eKait4k9hpdtqTM1zrsgYT4fjWTHE6zBGJr/Qk77WFKZQrGCorIIPZf000cewj
2tXoJ66sXTRFbeL9uw1BhPto+r3QBX6SlhiauDtk8mnwhbx3VDi7NJHe9gkjmmgwJx3GLvZFOOWX
UCm+CwYqgzzNJ8qbvuO2TpKPNw+CtMHDAIeA+Y4jKp5THcBWXY1dPaU+V530fu+p6negLikNQomP
DFO91DKZz9zH2t01Sk0wEQF7K0jcSIxJFEoYFQtB1DyT3rXV4iq16f07YLuo4E7qfllwETBc24Is
SckoiBFWdY8mT//aaN/Ox5DtcRoOupW5jhmG6mrmzT1WgB4T7Fbemgy3G6X2Ax3CnNEsyNoZM3tO
bDXWjJB67QiBm+3PUHvchSa22j7Tbt05gBDjqiUdtvBeiG8BlQ106TkApV1P4n1SoiwvStDxcB76
LaeM1KH/ifh2U1LPbEZjEbNVc5wXIgJbGngt64ILV8DV5d9Ceciutnakcnziq/9Xh/JekKSFt0Ay
yTXv5uMJwyH+omIXg6nXPTqt63Libh3B3fupFyVAAvy5welV8XD5KS265BwyDhSubIYok30C3y+G
QOSETn58PjEWP/cGq+8yeGjSwME9zbRZFy0e5cCYBtWXY3oXvGoWAD9BS76SOflcAs4TbWdcUXGz
KWO3/EcNOYWodkERivTgLx+UA/Ni7hu9WgTZbzhd5V7nvqYEmRwnpzPbozTQlYXADOgs2YrOpnVj
MUURX9E/HGlOfAg0CoGdtkmJoukO4zPSgqZ9nlqQxwuqeEnZXL9A71mczdKqE2LMQssfcK6IMCoO
FEnQHRbrhMMGmrVPc/Ita3aQIYimTZ0X03JQK86QA0csKPHasEUW2ZcIi2/LjxX1+jVF4pLfOudn
DU+7tlpEELTljGXpNrzfW02gyPNjDrwJqgnjLqSeI350jADgnhWSOEa8DrGq0MaI1iLgM4F/ifBH
IW9AWToe1Pg7sudyZSH/SomVytSo0jatdda+VEWuNZMbFDyI8LN+rKtIbtCr5r7KYE6UIhFjkixT
KG1BfMtfYkib21ENLF8jhjdmbVO7YsSJfHDrKWCl870iwTHjbTMSgJ8LNosAjFEQLoLuUvuFKGMh
ek3V29aBQei2EzqcnpRguSEAjnp7KENIPt4l+b/sd13cBhdAsLa+tX6W9nThicxdi/R04bVoiNkp
ieC/gDgL2Whb9iEFN+r+hHzs5MmbG68CtJRPta8rAGqlX5Xq4Fv8nIf6+2OcHuWN+9mOJ9QKyzu2
lCGXruotLnPY6q6Br+JOq7h1okaYz8tL6Y+lmo6WeWmH7Vn28y16CdL0ZXSxWE2MGCgWwpLGZ5f9
h7lmoGYHX2Nr2Chnssd8o9SC9qzy06aFPhZwNLN0wR9PveuEqyu8et7f9Y8NTw6URh8tMThEaU0N
nEo2nwg57RTNZzKwAWAylx9i3DOOH5v3ui7fEPJz1852OIb03VareGamO2dEZXjQo7khX7SxWoxy
zdj89rvCf/iJzYdwpRrLq+O8eWTSZGNqQXOTeB0wxALWDtuNhoA9dK8m8vTt9gPOixAbSydH2CpK
sdGe2OdEs+2GMXnpsxWpYLeIG5FLREh21Uiz5aHSFy5PcXdFphB7lhqkfe6fGVPgUq67vHfbeMxn
Ff6Kt5H3THaZr/n1eUh/Pk0d1yj/y9jrkqeMHsueqqggw7uBhaY4qyOlblezf88ccsgSKxGGb3cB
z4AjVx2wmasEcXOzlSzmV2VS+dsNsIBWl9nvWxUTIKPMM+QZmqqG926aYYEnhs37a5+Tcffjobwo
Kt3YT32FFHlvkbzHfO7YtiVeUHI0Yb2EpNMIoK+pyniR1hY6LdjqLoD8UBSSaBshjNMfq2svG7Z6
IIqXzcfgyXljfP5bvagctiGB8Y8AhQ/5ZWaxMsvz6Xr+s7TScsbI/6sEjY20ZsiMfwAzp6CFhO1r
2BUmYYkzM+FKds7ay3Ds6jEJ71Ad41R6xtBINBjBOhvTkloidc+GBGbe8VKt84/Mjktu3KUGj7fX
Qo6BcWZoo2bpRkXli8R96Exyy95lAuDtUnkMn3/XmKZHUoPr56B4Lf1gnPbOftiGiyWAM/rdnFgt
xQAAQV2CEimMlY2YWGPNJDybY915rsCIr8aQgNo9tL6exEeWxXKPyzaeTvnF64x/DSY953kDKDeU
R2GoxtW6Zj4uQuDIpWT5SzlRZxVB97wsD+GaZmmPneE+moNV1r6ySly5U/uH29sZmqWVe5lXbTgb
bjbqKb2qA4fX7/dVTi96stlmzUcCvoXx5PvIfaNLvgSuL9FptNQP68Qsrfz7I3r/L3ySJr9jyxIa
1ri2lEq4S7OBZReov6HTo0jyFHsV+PnrMklMdlIWnHSKMRlt9qEnZH7+XLtkzBLVWiX0Vf48cBwZ
bCnDVucNFOiUQKSmIbXb7Iwap3OUYLtqrrLbKm3YeSxN+FIdytOtyWjuPEZkwsplY1fXt6u6Jw0Y
d2xHOKPFdp435BPjaqCtfBsGWcHoM6/jifTCfGq64FsnqwrwfKWXEob5l6tzECgp81VgQDxxkGxe
7MgtXv/FG+cAtuvqPlSfA58VUVsLXKRNf5MaPRoGTkE89ffLeMx7tIki+L2wYIX+bQEj+Xf7phhx
kbvstIq01svenEbdjS4r4GxuUJxpd+szAtLkxmVGTVFLvX155s7S+egFcnmB7OS1oqvvxRW4rk3E
NG5mYMIEqOTqmdRRzwwSgevWzISOAF3M/biTGfrf1Xz+eECzJaKiY4mltoGkbq1Q9vngUXRz2qFx
niqV40/Pyf1SnQChaQ2VGqGG3V/3Y15eIo/HmGp3wx+yjuUbQNxheXwlH9OpCpq7u//LXdcLZT+Z
m0KyD99k7DDZSpcswnneM80StZOfZ0VwlxYvgWk0owldgjs3mM+SVk6fg1voQYswuP9u1brgW2L/
Q5YzUgvIn6JskASistMeDKJNfELBeVRyIajq3biLwio2ncIyH7mpoXmrvmT2jOtMtU4eQAoq+VM7
/4VdAx78Hmj9J+R+32hXHfBR0v1hca3S7UzwW43IjoD6CUKycOYC9lz4hkqOwM9nqlpph2CMfVfF
0oXAzXe1BVeXRUkTPjI3SFPqlSQNO+BvG1khJqfn8P+7vULLkhPhmM/Ko+q+8xBFx452/r06zzbX
YIZ87ETiLACzoKGcDvkCW2/8Nlgi9bzagdB1klidQuodCxY62c8SP9Jy2sY3o/hNqs5wOu71fJo0
3waVJiezZb0T9jzARBwViiI2i99M+LzPmt04Tcyxz65S+cpb1bUfroefn5GZEsz5NmP15DmnrpBJ
pG77VpnHODd8zfWBu85Eqml8hzDkNUUgGKXcIAuGRlEOZoeoOItqsIVDfhrZilo0FicVHLJjKsGH
GF2rQ1wBy50ettzr9KVOGbN2w9Z2rXMa0pSmj1B64qcMqlXNZveDc6Ze0TZwjNX1Ip24V7NXMFJp
d5AQL0XHJ0mfdfmx5FGGwYjIGTlCWlRclSe2HQxG2ZHosakEIcS2xbeMoVNys1NgbJdh9AGadXWR
HkKaHNpligb538/+QzTAEXEWta6cZwBMGMEkh2XnjTGTC8OoOsDUVNI/jkodktpkYrSDODcXrogF
dRgaVfvi/09lhQUzIyznncupQo/V2aWVn+jlqMQRiyfDpg9VAr7mQdRh1mGmuLvcGbiAmB2wG9mj
Ib5h4I7MBj10dHL9eNhvQxTfAs8MUb4w5A0wIROeFzH0xy5jk5maexOQu2Lqw8uK7ANTrcVF9zzx
3PNp/xu5Ut0MTEDcqkcmuZfD1/knuN/r3YPS3elhvhZoiTzIlMN65vnj2x0hsbcFpQEUKcu0VjSb
femHMIqocUuWITNSTfaDf5q9Dh82jz+6ODfF6rgAhVwJNPD/hfhYP4CR9q4ODxUpH8d9nZiZjnlL
p3NxKtuSazjwfg4+Hc36amq+nPI2TQaRhRdikT1KNl7RDpPdLLY6qg94idQUA4Pi4F72J5GsXMDB
Jh12PwfBTNRfbdT5/wm6GP5IhI0dpEFsSbtIAk6GqfP1WWdD0qOTHLNJOqEXR+zv9ul0XD/9t6/M
SB9kh1q9u4UiVIML/9JyrvEjPrYF9560HNc4VnngpmOQm6PjZ25X87ifLQ2z06jQjXmLX0jx+vjC
WakRFYh51PMFZyECTXAS8IjmK9AopGj1X2g05u2rwQdWLJrLTW0jukDdF5HBUyzbSJ+el5TykREf
sIraigFlFF5v7ULT3ud8BHpjrNhOEjJt3utFUwzd0g7QIRXTAlHnUJPNLf1TiZjF5Sg4wb1eC2uy
3Ql1o6S4PR5xmxgpTCfmWB7D2yWxrVLPLtR+tU99Vh3kS9WTAXCjq7TF685HlBlvUp0EuQrUzrC0
/2KD1ahXYFDV44FcCgwa/qp1zc00jlFBC0vsAfZKl8V642OJnzHr4QForSV5ZvimZiw77ZGCysm8
JQtv68+7x649cMeiRDqQ1f3eX+iWlBI5gzHN04sv/zpmqMgk4S/neqb+93uqF2KaNMpalDUbXCCa
q81J/p15vRQrRCBThYAthGS6uYv+dG4LKe9Ad7Jd5zqKcVKgDNWy77zXHEFwILOpSz9Loy1Q813Y
YkUZ14TMHL4hutIlnf+liZYcoETuSZEVQSxLRBYDUomGH9F3OEtWwWh4QkNg9hF5S5fnVRTi9OUU
ZltiR+5Ddk3qO/T8eI7zrIPnEzZuCOpZPICeh5I3RvYfS5bJvqtiX+Oo86aMEl/ujgkXFfm0b50F
65zFkMEpalONfNZsvDlCN1PQmvHr3/5qKqjOBt8euGQtNZGHRQLO9AzhfVNovLcBeg6oelkykeOs
JlkW2qBvUmjW97PFrOgCrP++EF1zKEBbRK8thGshPZu5SzGQBIjnSeigYEVv74h7/OkLOnBY3EDG
it2/UMq98GGZUMm669tsVbtyah0fRJCjtYUcP9Nw251Esr1qyWrmEnKRaYIKdOXXaNnXeKlcnF2W
Sd/5tqkEzpiWn0A0e7lowqrj3ErMtjYK/e01og21dWQ1WAM7IBsPOjiZXL6+nJ7rMJTpe6PkF1K3
PhCjw6hoYlt0oeznNZf+IefTEydO8XFLDzt0hF1F53GHOZOdqjvmPqZzBKoE6lZt3+rpRLLMP94d
CAWgv5hoat/PY1AmMdnP33vNQWsle1bLs9M3fCRWPyYmv4KfwvEw3iTSkchpv44du0ySCFISzv1Y
6SV9QkQo/2j9CrEiDmq2DTquR/iYgwFkDUTlzamu617SoiJ1fnecz+rfUf24ekE//zDa8QKrIG50
B/eeWhDD9sCy1iX9VCgvxrTWVZC67pxz+dK2nlVUTxtcDTqVCBhIi44ycwSKIlAKo/3x9pIR4cTq
khovYMKFDkKXjl2h7B185uFsOxWjQ/HE03P1c1jbaLGHNg64uky9L9odckzxqR/OImVjY1MV2gdx
69bRFSUNG37acNkJh1Czs2zuXzjFZyebGxNpyk76kZoujEHD6AR1d4khO0pwTOgcljcZe5LPbw12
s0/HJ3dOeFKw0i/WSyZXzvZ2UO5FGDMka8PscLWCibDd4rap3i8Bfiajasc6rc3ZvgTw1DG10J7y
yKquFW7MpjkPaDD8OnkqLY+A6q4UWuVZimbRF35jIOT9/IPVWdWQOItfYabzhislpPXqcjxePES6
tKyi+S5d2Z/Kdhod8vd6upbsXneYM5pE/vi+0cBqupiTl2vbOtvczKljblj74/Nyf1Exx/IgtHNU
X0DGjywj6Mb5Di+Vrw2ELN5haeY4KF/mSTiWGZU0Qi4mcHhRuk1DfpkJ7O5Wyc7o4u1EJGtn7v76
9KzHpp+Hd5eRaxWnwLUrLIzOIB1UMSoKv4OJ0fxuZQn6AYhdOLISUXIVPvSGRqvqr3Xqo4I00KAF
41iy2uR8avSOFC6hBMLIooRk+RrIfCq06EvoV9FqW3pCAkXu1LvJlEWenoO5lVXG2q4D+pONeIsU
eOFvXv7tqNgx5noiikF8xjw5xGobgQJJubxokhEbUe7p3Vz2uyBsGFlXKiMMnPTTwtTKQ18Dpf/6
j8MEeHwOy8Nm1dZfvrCvy2v/S6hEbtH6ftbCSZuAFedO5TTfwIJnw0cgeISdAcDWv5MQqDzWHDjS
Z6pU2YgREaHxULqyUW42U8IyOphkbsP8mnpkZb5r4RmKB29TREIuKuuzTD0oUrWSUyNa8nv/UMh/
MDVijKnrz6zsmFZ72+sPPxDcO+vnGViPTjrLD0AjvxwD6RsuRf4EIQdI0qD599tDEEJb57vbRlL/
HFgEYeZixAj2kpGnOMrQ+JLP6znOye6UK5nD3zwJTT3AtPudzIUB3yt6JtiVtp5zE84Oy6xHOnGV
BI2PtvQqo8/a/FW6UysbbugFCJf6mFOJBR/MN2CI+I8am+4T6PMnFnMySz2W4Z5OBZZwZK9YP6TY
77pUcAoEvXlymNB6T9Oo2GwNfKcNMQFTMCozYs3jQH1dl9PqcGA+Fe80EV87lvEa/eHWTPD6BFdt
oHW/gEu92WwB74QLn8YFEPz5XBc9DhH+eILkhk3d2tbBu28lcUSnW1gTtyac2y3T7dxXeAuhdtwh
nMFBFa8fSUhn0QvmAb3j5LnPiRDRrC5I3nmGbfhmkgmYU6zrhvy10PTLtLOrAbODhU5rgHkuJgTj
F0WPfljw6JMK9WPurwXX1zXrVhiUtY32je42VzmA4kcZDofV6pbl3ALV2c7m03gXPP7bE7wvNO8X
+qiQzEDtDU93oYmoGJC65OnpgxEVCYqczWWqSg1iffn8zZuENcF73pWcF4aX9VVkMRcHXmgIuXHS
y05jLdhZYK7X9dezLi3fNgbfZ+3lvUdc5EPdINz8XJiVkYLKChTFvjP4W0UD5fVgOKL4KwLuJ1Rn
fgN+YjIcujfyg1Det8O0M+gFD7G6yHd1OcDep77k8P3UyWNQsLTgsSQ0qUJRC/ogZ2bBh7fn7mcC
l4/Og4FqgqVnxtoQaGEGez7ymY8QXJO51ocs/RKHz96BJgbgC8CxOjSWA/keSkai/ayO4kRPbU1y
E3+MwBRPn7aDoDkeEpZI4MW/tamNS3W2S6DTHz7EerPt5Xm/Co6LpAJcEZazGelVOSKMBk75xSqE
tw1u0QIgwDfAiyElX1KDqolSN4GyumIoIx9YjRMUl2+4lA/mZOFgWg9K37vtToL70iGBzlnibdVL
0zbF2XYcQPJzjqExDShgWCSpp9yiRTLgul+Kc4cC9EVaN1LylracYtfVzbImqmQjlHEDU4Pzpxxk
YmJGEBZIcIkQ8FXZ1VYQqHgRubRtUIUj6RCeSCRIfscLNDk2v5U3MUgBb0rA3JMRUeiuntYa8s7B
i7f2K8GgMnsEnlJ9btNjA6aXXHcFz1OYoeVXGdd+iY26Ug9r89mQQaPLcqBBUOhtFCWx1MLMKEdV
wtFTzzwltRBB6BGuPLdMCXDDDba7vZESYIerGRN1oE3almbYXcTcEPYHBHztNgG2ZG/EfHLRcNCk
hK6Pdu0WIl6khhSWAIQlHrdY2VhO/Ou23DQdslixEIoUy1tgHwJGyIokUr/rA9e89reqFmSTiyDe
sOVi0n+7xLkCjDw+0B5QV3yZMvYmfOQais21+emUEew++uK9muWVMWPKrpaGe9tMNSbK7bSrtvCG
Kf1xoMVyaN+YuBj2oWEOWb5VjKtTNcmfmAaWE+0gpc/RdVPvBeVXblproQPFh2FzvsFF9IGGuhdo
XqTzHK51Fwq9myRfPjKul8Vgu/8fwkO/Ttt/1hO2P7aG5FonLMhf7WEIj30EqUazTnmHGaq+kjOl
GDpf1TN9Zl3yy3fsdx4RkVMOJ4lSfs2SnBH2fO9P0hJkaO/0LQiaPpOpUWWdxueOpSMOJq+nY3Mi
D39HBP5tDhYgVAvgKKeWFUyMOo1uzgu9OALac9oHgLbIwVTEppjXrsGCdMNEvIFiNgKnCUyoYEam
BdEIfuCrHi7EPjG1WTHqQz1jMAOfxN0cNlmttGm9oYuWyZ0wqAZ5eppB35vYCbNQ1xTz/gUfhz7m
LL12V6vX6jLja93LQy8nyDes+5ulu1DeLOxjxB0bZyXJsaRnQANDex8aPD/FrP4xFqMDl81sa/4x
zgbncH2yyGYlwypLJs0DN/97kTi3woU/5HK2uJgXaMlJ3ENaVi4f8evdafJPCU4A9/WrHZ9dg3Hq
5Ntnc6MVKP7ql/kJ7rxRXTEvyAbqUNIdgT8NVw2tUxNYd8VNbmExUL3JWjXj+k4I9Pzz9kbInR+n
RKDK4utnxd/1EasyZktitWULHoobNaBWgG95iBW7/m4zrT19dIdvXoBDw9ycYCxuZKN2ZAmXGraX
sm1VNhNdhL8S/ycBk1OJATr5Bugo9f1aDTfCgAH6QPlLJjDPoh4AxcADO/4yzycXhyImzU1qffHN
GDOfKFNp6MSs2IJX7e13Ut+NHak1kMKi4MqjJuIHEjUNQZ6m1VAZOwibAOxIEJtT8uwqlwxWL4aw
zaz98AvBhscROLQc/oQdD3olp+1b8si5TQwRE1hz/AYq6laul86xg6euRu7AF9zbL4wrUzoz43G9
8oooj3Tf2bKBZ3ZDfEOyTPB6DCKIHQrmykdlETx97/NMlknoWaEMvF/i4XHS4YVIOQYBAO2Hk04c
HA5dz0Uft++fxkozFnBSCVQ55e9UFqluUX/m1pHXEs3uVKa0AjLR1koWQjzxLQmAS3HGe1Ob40wo
tk36I7Kfea5OovXQBCP/O4NeqDQFyFxpDMEACexKsjr9wWyNDRYURg9PTTSr44/FGlOqTIsyw3DW
n2Hv7cw0PSXR4+mxFicgKwRfktgcJ5Fr7NmKL92mxuRvLMeQeWEpyn20BIeaI1GazN0eN0vtGGqE
dXGe7nmVPvDulB6/FsAVmV+N+7ua+Yl3BDppkIce/Tl/428PXgRhXK741NAGIzdFhwi3tCTSLNV9
G8PWzJjmIN+0d6bsToGuMmiBljs0ZwRbsrdr06N6lvjsMkXQnfzyJSsIZMElGpjfaKHRy8mHFJO1
uzqa9aRN/eP/eQR5+wfyvehTa9hjXIMC62PFn/QofaEM4N3vqARAodxcGiwtNsn8qnVtoVWquctU
9OSIA6LgzbDyE/7B+R+MgwN14lW8S7wjrROT5m58l92YSS2NA4f2KsCmw0Sdz0Bxay9ejfC9/7p6
4+Y4qw9DOy5Uz0s14jGIJYSnsTvEMyF6THD3G8S23JMYkKahEtSU3ssbCfIIrKS80buPZb8gu36W
KEinKLV0PsPQ//smtIffH0ohaZr2FXRexpF75MHIg067NkTuzGlfVhrIaGivmm1/URFZ+OGwBqZT
ewARnI/2mDVprBy+lGtKhI36nBn019Gip8QZb/Zz4iWGK2G6Z+FPwTKmxYmjEpEomEr9JIUKkC37
TBps79qN4hzEsJLXgrIXtFv94lH2/qvQkxvIdtW/+5UhhGL0qCAMyN8mes1q5LGoT3dGoKlwjEzA
cfHuffOlVEISC/Ie179PGqnTYepMTVXK+N0EGs6wTeFWx9DYpF90BRSXFtFPF0HhtimSoxsWN2wy
8ubGtrjFgs6mVJlcdeTp5iDRZZSPP5vgFiadaGDsr/JEAuMY6q2MGJR9vcXTGMlZzKrAV7x9Z4dA
5ZIHvFGgrumTAQcwjXTXZ0Fv4N8qINGOCXOBDETNd3Nmb8exY8i4V0TDrD3yfmQwEAcQMFCd1AH6
ILDZPVuLiNhelj3yg9psyGYF5IzCvGyLt5iRWBX6x/nDzFsdfCGdiAX2MuUW80OoOR8urzNggnsS
C3OsPcdX+EtZ54rqQSuqFjJ6ICr15ZylBauXaaI3oh5w0seqplM0WK9Hxu+5c7Tf6W4yNfySva/X
38Sy7QHrrBE3c43iWPofu1fI20dwQTVoAISvmkaY+t4Dnj45d0njSd+hKSG84ff1L5SlYR7biryu
eqnyTOxF7IW0sVE5xNCmTETijcffVdrVUY1pgsCxOyOBU+yZINa8WRtoSWl+dCFMf+UMi4LiVpF8
EKDzF5uC/eDKHFCGPcadvYPn0xjbdo7wnt9ektHH5NrtXFKnjbr+pZcv4xU6R5eghxf8cz1k+FEB
zqLMPLdgzK2YLpAwln2q19zbqylwj02OT7oe/GNpzufkMx1kCobgC3E5d1VPgbe/mOrS+4dJk3xu
IVViuwy7MsuE8I3aZDcCABkgdT7JM+pZXLAl+ZQ7SzGMWll/G0PVCAwkKLmvkz2mgaHed7duObmH
AHF131H84WOhUhUPV5l7/Z2K+rMtxZ7ajTqWyNe09Jag1lYxdJRsNVTiI0I3XYDJWeoFfPZnJnqH
2/8WAW0o0HiE6SuRUBkenUZQD/CIyqGpTwOFDTxkrTM4urHYBcpTM/Z8rrfS0EB0sbOptEldbgqA
Mu8rD8t1d3McBPard6ATDpltQjI1p2qsf0wjMrwiUlW1bz5/Gmcsa4+tYiOqLYcix6iVvZNjJg86
rEz6B042NvKhaMLkOVhYq0uvcNKECdaQ6byAhcnvn/F/goTxB4cVE/FqWxOZy9YSsvq2bruCN1Yk
gCVRA/QWom6STxsPokbVwxYfa+4Mn86yKIq5B//1lBAQKbHI6T78Ar6w5Oho8+0zdCK/5r1YD9e0
ahAzXDyp+XjdxLu/J7d/o50Gk9KWvfWKPyaNIZHjij6Xms0Gf6UhaTieSUGBoEjAmzJPmmee7xGg
qwv8lXOyX1wn5Zdk/Vl2cJNhVFDgkrRUlFJQeg8R8hr9rwZb1QkTxmAZ+l3dZ6D7ValmfCE5akU6
kMQOZ8/wf9zQF3bOYGGmFinbV/mi83ytd0sXswrsy5Z91IrQQE6J1YA0C8Ph4QGboWpo1BOjJzBh
5Xr91+lb3Qaiidv20PcMGzROnoS50U6U99iMRCKphsTpF+RRrAPQwcO8fWcOs2rZ7MqTQ2NlKfKc
3u2ia9ffozwvpeAGAdRLRNncMzQd+wD92il/yqjttRhi+dykVgYY0zbuGb39BaftsPvk58SrEg2q
OvBSa+xiimhZZmcu1EF9m1gopC0ouF3J1LuMC8uVBeZ70DM0IvnCTusnt6cJ9pSb/99L1ZRvX9SS
ARKHrC2jN/dT8gIbgs6VdIm5aIeRzqMlkcgS1ageAySZB4DQ/4mdFSdtXcb4COg9rTusyuYgR2Aj
dSPnuqLhXFV+Ry8KP7gniMRoFuvDa2ym3MGrUSRP1GaDJrPAOftfaYyGPo37zitx69MpO5uR8T21
9oDglIcLgtW9BdmMdESyydd1rU1QWUze9IVQicbd6V7E0vY16qRrfiX/LUeS5E5qRwtZ5YBT3Hv6
KPYy8wzsMRHpsrwACslCN6VGwwwzoKKvPWrpDkGf1fqywF7oWxC5wnjw6m6bUKCKtF67XpOys1k8
grUMa/RAI/8sOz9zs8/RaBg1FwBeRkbIle68c0F5bTh4c2E7glan+psVOYaJmQ0Sn57Y2+BHgJ3U
mAiQJGtLAZ5BLo35rx1sJhPPivpewndoFixAOhyLzfK5Y+GyYT/ThK6BHqOv7IDzkvc9lvVL+MBG
0/8S6YXrGaEmqFIYUcAlxlAsS0VYhgyns4VfUrtlFpnCxu8DzLaH6aZUSw9hluZWn4cMFhAtXX/T
me4ul+yY3ge6MZwXerx9yKs0nU4JNf/NBP2A4bILBsepVDnx48eOhA23QqGLXetmu05oDkqi8uvL
aN/THc5r36LL4rTPWLGKS+zeVecfE9SZU14NdBppB1IgaE6TzT4ruPUc97rolJ5FoRYnSnQKbLkR
JKxJ/P5un+0ffWngmNtuAF0QZHj9VH/H7/gJEK7zTAFcoIj9MSYKkw5NuhdlibV4MFalg6gnZwM9
unGkzKPcc6+e+vSpTXDUX8b3lzwy7mrc4aY3Tjz/fC8VVO8e68BmGtbELopUuQouhDyBjFdyvjDK
aMZVdeRA1YrK93zwjUPqW0ZZThAK4M+hVhtXKrM6Aht8BqMRzxrjjnlbNAaqzlUAYCZpqfNJ/LmU
f0dWB1kX3TfAeE2evJvQ47AqZgSdb54tk8swT//IxFgSLU6gYXtI/35gcMYyix5fKvqJUfdHFxgd
V1aawHlALj9coPELEDvQ92H/CJ8uZJ2ePcrA9yQg+wma7zTqBVzuDoqlkAox6DnLj4COswVdy2wQ
v9izeJNwiGgqdDDVUfHqSL0fBOOiEtOu8hBy5BG+/BzJhvtVdWXUKXPY/mhCpGkBDLDodDjvMyFr
rDwd/iW4RnOB11EtyQu8Gcy76xjyXJpBKh4SK1jSdElxjcceTrKlqreOgAsrDTdleGU9otWFPeT7
V61FQBXh8u4feCQJNf1IwmgE814uvIfjvKNODbCJmzSC8s6RersNH9ou2C7GCvBY5BjznhaP3X1P
ZfNdS1yRjd9DTXepUBJiAj/YghFOu9/Soo2ppQXls00hlygB3rbf3oFzhRJz5PWRQ/8cJrJw0oL+
HmviHfZFOVpyoyGosDa6ImjpIWU1QWCOlFkrbYUMsv3L0I09S3LECXheNy72r3Igl2uTDfP8XFJV
qS/A1SRAo/WhxsK4FQ28TqqoFoHwugyk/blSvICRnmWiti/fTcfSXCzlLKpl1uVgkyYDRzc/TzWi
LpY7R6nIOFmOdK73rXvC8NriJDKLKB8IeRBnSCx+saADym2Js78z9O2K+mrvrSM2IbThf852dYdV
5hrVzyxTMnB/NUkEDvgEueNUGmDAgzDHVnb5fkwMlwMWh8S2l0qo+oZFI0/OGdG83BK1FckZS2C5
jYT5uFEJe64pCRRmm7QsmCoReb+jAYuHu59lSDFwgwSJQ6zZ0Y8AlR9j4bhKLTTlZxVcPIt77EYJ
jj5YFKsTYGbgvVp8Va/7jIG7M7eMa8rydCrOEvwKhnUm3pkERX6jFhGCo9ZSPjB2QfHVanNLJHEt
eOVQoRXT2ebqGo7hIbPZF6vHZ2ziGEl7xVoMpO1khqfVs0dZUcIQp3tI2Yf9QwWSre949l8wRPIA
hDtiT13F2p1uItE376OC3j/beXJZ2IeY+hcnN3Yh65sZSyFIJIba+Z6CpRTeXrohC9H+PTrvi48D
n94vLqndkG9yN8Cstdb8EO58oe4l7p5egCuK3RNH21nA5ckylpUY5cV1REWSqhKKNWSGoR7guZCc
TB/prJvXAx+wOl0pcBTxFFVF46MZNCAz0rmrZ3fxPzyxwUi6b2cAciCD1ETbB3/ueyMrVYVf4Oh5
GLqiLzJQZK76VNNXEIfSucqtmqwe01c6cv0gRlFNrjqYvUBIREMxkzAzAoBtnMV28uBw4MAEB0zZ
WlGbknj27wy2urI51rNxt8CqWGzRjhAPk253bkCc+MZsL0h6zZoLEo7SUhNO4c4gE9WgfoXwoTk7
wuTvzUpb9ZJFAhj8Wlq38hngpmAtT329lDiOHcCjHZrjgh99ndDYZgeFaWxaJQWd+UGnCHVzZcLF
TRSZYxVMmwBm4eAdWCYcn0TlIcYIcmsx0LSqYn5dAbZHUXKNNmGAc8KXvUxxkTsKIpxlcu1ydDqJ
g3pt6Hg7X0wgbaxvqdJMLS8Wh+rl26p8zb8dBAOEUNbJdD2bdyXo/gIyQuwwTPBQfhG7J1LI0tWm
IiP/cx5HaRZKqXlx0x5X1y/zdT6LwWOA/QwUeuVoa7zZI5I+oP3jmJo3kjc0RSYsMacrFJ5APoNj
raBrto1UWbazQslteC4ssXlidZfsVlth5fVdgccMXVwDF9DIuSkFTJynM4hd72XQg0tAS5l5cEJr
pSjlCxnm1vquKecRg/OW9tToNFZnqaJq2JMmcX2OVaf+flKAX3SbnzlGzGTxMG1+AnelujjOtEGZ
XV6xZLeS4pn88ZpSquJzfZN89rcLnPtSS8qCK80ZZZNATihw2akkrSyzk1RdKgAoIhN1dakcNlot
oLhglLto6QhMslq1gcmCzpzNpN1KhpCXWnxXdlgmC9KfjlFdx9VgbA1sMDt9YN8v4NK+fnvtW2qs
LRnwFeSbCZq48aenW9m1AG0+cNI37hlV73UAPV5hbgxhQxzbOsNT1DebJmX+UfSINML3P97ep3KR
4oxCIypXxXIA9FsU5pCiiVYXJ0AwcGKMnXyZP30YlWlVYVx5nDYUTIoeUWzb+qHiavp1hyC4ZWWe
DmAF1oqfSAqzY/PK7vqKYdJS1hm1llTq/n66j7X9dNtirQPjUMbrA/4p0/d9CYACR1LwGdlbf8wx
evixUKvrUeOcdOUeUOvS1qANeWoTnGSckAG/OnZ2liHAPVfhAYmBRxd4TqQrwHdsInorHsO+cFL1
2ndCY6X3RbiZ2rlL7bY0RGw235s4yf0AoQWYB5yrVPmPq5RFGPbLsKCrFIEiGrMaLs+vln2U49Wb
m7TniIvXldzsN4tLcNy8GURCSLOV6AhZXiM7Sz9/Z7Vhugg9nK6GBZ0iC4/lYTtUIbRx0V8241L7
huysjmYEdNGKDOvdhChC/FO7hgaJIwu9aRh/bLz5ldYWjTpYNxPo8K8Qjjido8fh21ecFF+bvRqb
abCPr+KDLNRSRfDXMnJkb5sdU2HF8Q2L2zC+c2CqPQ58lL18X1VogunjlmRmcG521EzmpHxNVCpN
yxdexRxgQ/Y/tJyrGJIwpBbD1UtHLDvr9h6+EJeXcX9lfRNhlJm8zriNK4WpYosLuemd3sfq1DrH
zSHf3UCzgEsLKVjPAqmsLtMYEuQfF8CkBPNXjING5M65kA8DjmJ+XYF+2MOHz44zXNvHfEhSI2Ij
m2wGpuLTxZv6JvbphSkNlDTjuQN2S4yfZV+atHElaHx+BoiHFzasyIu4eNQ37uvxvLRQgu7xVcXy
qvCkEc8JWdsjweyL+sDkseKPsJil1Kk1rUifPt+9qtBrRj3KoXLL1HDrZOoLT53JIgRKkQcBmNA1
mqu+DJj8kDolD8WS67o2xKKdqnbnNIov8rWOknK9hFTtvEI1Ek2ale05f18ynoypjup74ulrrYK5
R6XKHsEFu1HorPtIY2MhoCvi4yksCwCbSKVJ+51OPKQFNDjPPeUdAnAosd03nARPZgSXSsV8GoQf
XL91LKSCK5j4GyIdM5SdxUl5lz+9foCef4B+8ROYKaFv4m3XALtyfFc8E9qytwaUXNk6OxXv66U5
3fNGRB+5mAcf0o0DcWwKe7jpN2Yjl8FwHp6fcat+ajIBq1SWFLwEK6Wi5d+h3rSKh6H8XxTKFZBo
EjiSJUJ0pKrMqCRdKSwyXvTLq9AMgBcLiMjiVFLZC5qQPM3SVnwdjjm+h9Yro4AQojGS6tA5Ag8B
ZNyiDFQT6Yxjc8w0AbcsJgko3Fz5xEksp0LTVZgqZgtY9Wh0nTm3i2BeLeIYINQCWgnvBnhleZI6
yYWTb2duBbNVIvsf5my/f0krepij5UJuUl5EAJ3ztIe1K8n0JYIqMLYHELh1gZ+93LMwwc0a9E97
wvt1D57P2CTnWcm2JIWvc8kQQGIXTdZAcN91KyOCxP0Ws0FTCNeOdLHqNS7F2PPss/ZoiFB/S0Qf
fr1dTpXAqNb/yHsqKrwwnKjwkFJJV4JxtsjL+smgpc5upP9GGMcvw0YHJJa5hWta9U+VByQQ9+/n
oQvAOrc2HkLasRfO1AkJk+ENxiTjSPTQPNdiJbOrOpafM7m8mtbCxYeZHrYeEsu7Ez0A7k1aLPW6
qPuHK6fe3ibtPLYeQ6jH+4+6lHNwKFRBlkLyotovjdt1DxxdkedVJSnc0OZM6+WZT+6xnZD6ZI/K
0CUVKu47fUTtV13RuQnNpmO45OyEeUDs0DSfo+R1PHj4/1hLIARhO5RbqMfx60fizO6rLpaLDRul
QFjdPqwqreHeCBlRWPH+XcXqqIM4XDvBX+lPacocQ3PbTpQtcbhwdaPmVLqBGtpliWGE+OyTm3Mb
v71//tI9Qs+/uKF9UiXLf1tg3OUfldMuzT9SlfEoqszxIfIJXP6A7BU0JOegM4ZRzlu3NAS8q7IS
9W/zkPnnMtqW+5atxiVCQuOdNfkHNCNKNi8rmMUUoiS2VY0jH8XDk2ZOOsJ2aOI/WGN+CL27M6UJ
MenjNkkOFwYUg0kRgDhDKE2ZbhfF21Q9CbcTi+vT/vl9dQfbv/PuyGwfF7ShHlqrZKYXoN+Yk01G
AEy6AsDK5EnfTeuYYMTzNP42RZHiyFe9V5XFmP9m4q02T98dNx8gyfZabjxFA5gqdNLox3YXwkbn
5TLNWBv9NzkUrhgc63WkE67gGLBfjXvUWpbSj22ft4ZydJNnJLerYKghWpRdps37CRsOjiNhYZxk
tzjCK4xfzuyGMTxVVao6H0Bkm9YwtToNy58PqfjXG+VlrubfVQsxE59vMzQk2L1K96tcZ2tBjGpg
+qCPJHOHDgluhCvko5J3lYBXhZg1geqGXOVSDooDfoMFLkuKYHoGkbUCc2/GNG9IeT3pOBJLePzD
b0M21NXpGW/CdoAkSwGvYceP/LMqGHWpV3LGrVeEGmSS1bXKL2P9vp3Y3WjAvZ5jp1NBn4IMNu38
ou8CiS9PYzxsOZU6Uh1gUP04tO9gwiwfUM71Vf3Xa0Mtf57bfXkv9LVhBDo+eD0xnQXTiejlGl5g
JZB3LAsxMZbrEWD7CuTxKmaT4bR5XDu8R/kNGLsyvsDmJ3frTt03sIJq+ypgk/Q5Lu/7dCtFYEsT
Rp5sJToroUjRi7qTvXlMXZ3n2N96jB4SLhXG+wz7K3TWHkW6z7p9VlyjBgxos3b4ajZ21+JOSxI/
tmS0tLDJnNFhkESMhFtXvOFwz8mOj6RXS9TrWfPe/1+CIhHFwB6olRNnijuWA10lsPe3Tx19qAC3
iz9EIgV7E5JAa4vyfnXf4YBXd3Ifb7LZJaGOccRB32RvsGms1iPKF3+RAIGPp1+wNE61VE/qTmQb
pl8EQs+yWjD5PIxK1HCbxlj2Qkew8qmtJKmlpZRt1xriWC47/nXKD6OBf2u4njUaszQuLk5+W46+
bFnl24tIUCMMzaEz9lYBDdj/c/tQUieuwRfehqluwn8b2MVWnt6Ijgh1DrL7o9BzVGo9ZGVcNCig
/URxGxj7R4wAHLOddcbj/dq+ikRRU5baYql2wwF30bj2k+q/2eWLW0CHePh+PQDmmxVxtmo5s0Ju
6hvZB9S6BYsw/UlJHFYr43n4GVyEvcqZ5vDFCztPpDQ8juesM5lN1jHHpc4RjduER46c2LWMCRiu
vr90wOn+GBtmXChyUzYpUwvEdHrmrP7ANyBzlCZ2dIZ220TqCe6fEmVLs23K0tkiy9bpF+Ng3hng
6BCGHZSYEiD9FKVs8e62Gb2JjQ/Ws1VR7zEFV3WxeW6nuBWHUU2OZDiyn8eein6PVAeWtC6wOp4Y
XsLDuG/+myBKtKlnaXvsTtGDSFeV9E8fEr9gwtwigX7r06i+yQx1hgJdm87AnO+W86BqmGw4pKTL
NnCPobhrAUDRy6uNZ1kolWHMpm+TJaxzfSZqSjkp/00CnGpX012b8n/6b3uXA8crnhmslyAIVsbW
EKRg7tZ370b+JIOG6z/2q7EOJTNOl+7FBtTX8QcJ1GYhs9YsIv4JgTVEFKG8sY6f9mKjbZFGLAYY
W2oFZL7zPL1PceQVGak2sqEtXn2Yg6QpeEo4DgoTav+ULHcvdwTxIhEXpSWcT3+lO5fbTMdJspRH
KKY8qkDN4PejxUM7S8U7Katm3QyWuID+HEIxLGKnTId670QqWNvpTKqJ/s7WnSvXEU9CPmvd8DCX
qMe5v4K65B4svmUhl3ObEFINb3nLZZDN05nC4i3fq7lBIiGGIvfBDCwrTSg3Sfn1eP8/Ie8iLSBd
LZ/Yu+HzgQct9GBLn9E4bxDLwSj6NXoN45cDfG7ijKZDXysb4dPgDEMJrZHT2pY+Ff97R9/1p1jy
VJ84hZtuezGpCJIeII6FRq3hgENrjNx6CiuCo1oryaX3Q5qK9vd9yc2/ryoHqqqVp8L6UP1rCL0n
1IqTrj5fit8bb2xQ8qZuHmm9m+KHdqpDmbdtI3B4cGvMB5z0muI1XGqGfsPcmKGXGIZ60Sw3Ydtg
t7gNWBTTvIg9C64zztLGvy9XgnhfE4MWSfAuxvyJKmAMaF4o7fRYqzwQwy6sjT7pv8SX9WnGVz5Y
yT1JylgF7UGZU82hx/A7Z/gVZUjEkFNfaS1wlbkDmKYdG0J2NaWBJnojv2EiRGvYRXhGcYf6AnC2
srtQFaUizuDNEyaPHFVFnZrM5YEt5SVMTd1H0y/i5UNn5ZOqOV6Tsb2xmfR6LYl9lRQYMukNhx++
nqs7NQHCWxbSbKNRKHyicnUq7UCAvgYLLNLLHJKHW0awB1U8/XfXLhy+/BvPlzynFfeGMeQppe9V
FceavCloK+o/9chKq5puxyyFmnCOTRG8zn3pJ9MeiEERa2nsJAULs5Ois9kpRUttOJLol6yMA/vF
e7lDvPAc/nBzTNc+Pi0uoUB1wFmNgTeEAvuKNRgGVU8ByN7dM3HcgYyKwJO2EQuaXdrJl7jpieF3
lFPBfXhmE+8Pykcz5asG3rJqfTo8c7EwshjbnoXiI8NLTiKgjPhRzSj66d/+GEomasvyEeZwA9pl
s7U6FA1haP3vFM9C9ipoF2BQoBCBZ0QBrSgTYd9vJnK4s9gEEx0OkfbyWjBSNikwr6lI6kCjs89D
GhLjecV72V2lIVvqt0EIrHxYcawJAV/tb9UZYtAwwx9cVSjqtuAP+7vOmXLM1ARsxeRAjWuLapmw
SqoqCLBx7BKo2OOhadY6Ad9t6omqQqLGAbZahriE59IyapvhBVgeakmZjBDebhIorpxkgFVMtXOO
0CrhvSAZtAxk6B4ABarc1KpTlNNXWF+YORM7WV75ngA0l5Qzj6bpQ3352I0oZjs2RVi9JIf7yWKL
JKPlvNWEKaxKImcmqQYeGn8hCI6jEn4EVw3foDXJ7Dc04BX4dUsT0/uQBZLwqB3OXwuJ+5YhOlYu
Z8gu3yHFc6B0rIr1Cdn5Se3zm2eD93/hbyZDmRaWqr6PlulNUDNgP7bvAyjtx+91yrhvUupxMS70
ZZreB+wB+BL7yyRf1H5m7jvdeM6bjJfLUJdA4g91mdiJJOEJF+NNrcsV+lLEsnS7MRV5+qEXwBYQ
j727M70TX040J9FLaWCT312nOooLPvKtZfdHEG/hUJW+CWCQHp1YpPMFSWRReKMVImuMtpwRBY2/
WfaQojOUWvbXM/8QPx0TJkqzBn2JSqlzn/rIN8FEolXcLEIJZ7N8Nx3PL9rFPwYMnScmXij3/7hE
t3kL6gIaSETiExmGlwpQxO3vnosYMo16D3mPGRxIoDgpqwWUiRAqWhC5cWYoMqP6BHmRQ6j/TCzh
K8V9uyuygFhXLFKTBVuimiWZhkGtd5e8vgqNXeY0bdUGV+Mm8MLdeZsBDgMzO4O83NIxFbwz8pWa
eBzTgM1FYGsDjekTPATw1We+1Ol0TtjfcNaVnq/Pakngt+mR9R5Vvz7+cBjSDfIlP+8HDpm5sydO
qPsJoBSnklxd2SIwi2VcWp47s39t16Uz4MkjpKuEA/fn246B4M3B6JziffrdDuA2tlb1RdI/Y/7a
9RJeXYRO967Y8ygMszrD0o64xOuB/Fo4H2dPF/4v1igVzLIc1v3mA9ZpkjjBOo0K4gsLVUsKkbhG
rAwrrYB04sogbgxXX/hT+IhbbAGtBlcfbMrF0MqYYjZI9ZmARWGfihd1fZ3Tx6STLeHhMQELW9A6
QPW0x2nrYhk5TTVMf1b9JPRiaW5yxl6HyHfrNHkLShINwUhlbk3nOz1l3lBPplZOEuw7Ukq4xnGe
TvSjOxyJGXzsDvKyaLrzXVMxwj2LKaONGsELx1ZaqAkXS18pydtlleQQc5B4fvrHhuDIhDcXJSSs
RbTe+WojXiz2aOYiaXlZIEvpEk3jc65eaAtQSp88B4mqTHCmgrbK1eBV+2ZjyT7urGjZVuNXpWYq
6tKyt5gav7RisvNlch7pgSeK/mGxT8+3m0nIzgDP7bpMkwIA2Ms7W24VJ3Bri8ffx3wkA4ySE69Q
B3ORWEViKEA05BHsYWxzq/QHCNo1qL4fYHJZ4b1jFb2jy1Qz7ishZS9ArVh6RUVL0bsQqtHa6tti
+B2bhsvwy53SRDnf5+4wrb5UxeMVx3MfisDSLdsUvQvxJbQ77Sstw7XJ7NInhpPyinzQIT3LbCYN
qp/+eGMztCxNVSdaB+Ve8kb7r2oFFmrDDABvCm8IrYdZ3K3V0V1idRWbxwdckSSsxQoBrgbqrQq1
XjKnkuw25HD1dNSLrSEmu5/t33v2NIjK/5wHH/rn9qmoYT0RJvAllUX50j72DXa6MOB8kiS/69il
XLR+/4jxxtm5qa55aw0xTcPrrHvjkYa7eDD6iUrsmtN+ZY3QbWkhUDUpMnTV0sqZLRSbWXm0SBks
iusIfFrgBD1PjiU4/rPbgXaxyJsByGbPKPoIP22V4ar8zaBmEzff9JOD7EDydt30zl5gSJHa7aY+
eAh82DUmPgqeVYa58Z/8SILX78Os8TqSqEQg+YI7kRmiTGa5BXXUBbAbyR9Fz53dbMIaRPcd5IbA
a1QXZPfvKQdn66wfKv3/y0JLeKduBdRpOZSBbWtdFuok7Uz/h66jKjbhJD6AFLlZLxSQCdCMZrTh
Z+kOqlvEdo/Lxy3Jk8a1pWCwJkPQccD5/3usJT465HDbOO2q4YapxBKoKL/IGoILtY1MzZKvxSdk
9yA7tQ8u6K+BF2b9W+8gL5QsfIh7s2ODNVLQHQTGCrXHUltdvrc54qw8XPoFpe6tXCBaKCz1xsWZ
tKqiBLV67FSfalW+t5pHHI6P5jVu4tL+qmxLzVcaOPrRTWJw/M7oEmMq6f4WIIs45RdrS7+ilL5C
vKKse22u/wskLVWSnkQaQq4aQ6I9qEsQZ0TrBrocguq0HT9NmzwInHDijCN+KCIaS1geUv3bPWZ/
YH8CT2jU7WpLhTi9jwK1g8BH+e+i5TIkFV76AxtPrR8mgVvVUJdxdOK1wvJwQtiETZiUcxLxyk9h
HVHtm8qIF+7qAwxUlu3/8m0U/UnV/8i1vmSX5Pjmfkb4n8IaaFgbF9ZGUqgvXFFlmXwmCv/r6TIb
tWMudysxNG6uva72HtJLHQjvgNxGeFQ8ROflc08WvPllehApOCipRiwp0CFCUBOI7QkIQIPQDQ48
HM0lZr/jzKp3ieiLFrv8JsfyeQ88SkTpKBpLh+GGAGcm+C5TmuGcBovI2hQCpjj0fC4Kyfm1Lanw
QsXyY3PDJP+P+1ZXAEAXZfZztb+g/pW06cyn8uBJjAeUhgARolLdd2sv5vCff9E9FuWI5jPNt94F
8qTb5ZaCyouDsjaNDFlQtxnAxgxFu9/sBPXzmLbnveDS0x0OAMZsJNCTRDGc90u9LNLeQJMT3cDK
dhYqgerLndzx6HzsiwT/oKYqARyi87BX3zWB8OVYgENeImD/3TVd3tk7fKX1hJjtfuCTu5GB+yBa
ygrQ5JygK8VtLx9MMkYl8DRwkNvap+AUeInbfFWbQE5Xy5PnBZMwTpyhhM77QrCEsRIMQpqW7hW1
JYtokF3Brnxf53oqsa8IAPJ6NWTG/uwyVjI5jnnAb6ubswJEnj7oq7uHQqqzzRgdS64Rt6eCocOr
earDvpKm99Oc8z3berhWel2PbC87QY3sD3y9rb0WgbEb1iApz+g+oo6aqR10mSU6V8jKUVJ64dt7
HXObcIeqm51UaYTCzwIvWXEZ7sa2iAKXGbP41ulq/R7jxr++NdGDdWlCBvxf89t3pi2JmTYJSmTC
EX/ohmfexLj4WqCfMwLclT44tWie+tl1KnpW8Joa6auNiMe/GT2co95QQ7XvpiHrfAahtr4rBGG3
srxMAEdSf8yC2utz5smqzM79Cvcv35m6l2WBlstmb90fsbEp8P0Nxtu2x7Z0gRGsE6ein8xfv6Ho
qMrWg4Qy57S0tDQDVa1vEKgSrXi5E5Oxpqu6JbHeHBg9D2rPSirJkMWe+qudXbJmvzVshkSMN+vP
SLsYAx3hxFsVBSMWmj4u8e6/lawAXHtZGmeMDR9BoQ0dE23uCfNDVQo0VNIRdfDNOJVbDRb/mwMH
EAQ1qa8BfrgEw0DgG83O9PXPV2UQC0O9CmWITnMwgYCLwpYK2OIq3cHBOPgx7BUJWYRpi4VShbhx
EksOhUFbcjCHtfWydq2RXoTb8ynTJV+IA2Qf5WtRa+e3IRTTJjudo8/Vu/9vMM9/o/6g4OcZlOaB
zZLbjfVZj0bWdFKGOS4Ze5Rz+e0scvlN+HFZn32LrU1teCZ447qe2BY4kuH1hVi/NMeBCdXWBj3e
oSPPBeXNlIun6DZhQpcoq8uEY1G47ovR1bBIsJMqUlStfCb2NhPGZV9goB4kXwAFg5XPmSLU+cQz
3lvEJDuNyff9YJpVB+Ave48gHr5wYz8YdbRsSSYGEhZq1Gra8cDC9Pyn1EccWZQ6CZ2LjXjMP7fN
03Fp8iUZFhKrfe75yZOsQAA2mno5+pm5DGxGe051cz9IfYINsuQhwqyQfH9G4swSCf1PbEydShK2
Q1x7eRhJJsTiEPUSfTRSk4kyPU6QlYdElfSWQsgJBn9Tz2dlrhF/Qdpf8jJAmg9TrSRPQTe3KGMq
qvWcCTnD/utbabi4p5wm/GxDMVPrBTOHCKHeTztqtCnXpSbCG4SSbLZobT+fnzLijG52uD0aNiI4
WYFH3ZQvdylcg1370T4dQ6dKEbxbBKcakBBrw3hZeM7XpQHRRvxfpPsdoD1U9ZTufzMgzWOnwLdf
qXsyXWfZMchX3ckx+doKIC5Tm5XY1vuHasi0LGuNbst8v26A9KyxzVEkK1EXLDCkh2UvMp4cQO8w
On+Fz3v/biTlqNFX9TZ24aD100RThFtyT35yJFoIzNyniJRb5Ap+sYU3Yqzu0E/xmCEPazJYUH/t
/SbZYdFEGo/Z7rQreR13ALK5Kw91rmiXZVxdT2AzkbI4YBY6xrFSc5/e+a6AbdRI9ErqoHBzshTk
RQh3On9phzZDAaEcDMkSodG/jc/7DRwtX9U6WbYlDGocWLLy0c3MUvMmsauG5cDIFBohAMYJFq5S
q4Woar5IjAcqJDzj+XwPGpHxD3bp5mfVDXdWMIHdSJ90O6M/tccD6OUc5NPYE+Ldqvt68IGpHt7y
PjjM7N6UehXvZR9i7UqG2551i6RfnJRpXgWR7QP2utof7V+XQphUWBg3Cfn7KE6+WtDlin7zef+H
241bpP73vK76g682tZyDSrj5G9wfkL8wZkHmGyj8x/kzSdcIM32LpMnFos5R2KeeSJtqmTqBDwvg
I2yZ7GfdfyMq27hYk/x/aqUqku7DhSBslB5OJzki4b5qhvhHoLEROFm5YxucLTe2Tb48zPrzq3iL
tjEQ9569Z69Tv+7+hDMTRTXYAPEgRBrIQX/+kKPFIhOVZaBWyDhCjaI0hZFQyOVPRIlOuMlAFqGz
GtdG0V3JMK7+rPyVlVF0ULdHsRj4g2tAHWCfUCyhzMBsW6HZr7xpoOoYnob9i8iyW53UtIvgywbI
XCpSRdHmb05RjkdsBDrTAJwnVkSaU4hyFl7f0xqg3GGDiop17S+QgBhgpdAhp3xFRXmRHDCtdxGe
LvRZlXBOndaBgyONK9DSPXA9b6dKUPVVEFvclvFUrdVvQzxYUjMGCxQW7lgnYZxrjnr9qzIz815N
GdCFi0pmoOXWnHNixRCg4ZLySkksGc8bPi2owSTUb2QqE3sDpcq0vqCC4JrO2INBA12JTxfdqRTM
ioU+v65UyJT/RPRXb0SbMiWarPZ2HUT1Sc3xft8SrX60zTghXCgBBUtzeRuFXric1VEihhNsZS6V
FuX/3+x5Qd1LR6/syJ3FBkPkSAKYCEWVWMVXly6nZY/H4uaRDewSgzxT+9R6hVwnfbUQdlHrPsnM
2o3ZvNDosgzVtaZN3Tayv8srwqeH3yh8Q4c18sY/eT9vOlcV6RFFjlquRmgRE8GJq7O9DgS2rEU9
Bhtn0xwHaPjJTVDSNypBHRyaGWZ6lgZS2BXvJSUvXfZgvlXF8WiT+eh2C5ebZH2nx6iibKJ/OWT2
ptbnaDNtvDFqEXDA0X7dKI8o6yN6VdBsN4/IeEkNrNBA7cJgYrW5ci9kRnUsTkwSNpvWP+K3NlVD
vP0rfFI7RNRTJgtgKIeeHkVTOxbWJcJ+vZZz8bJ6K23B75/izFxMVaohOEVCgMTqt+ZEzZgTcIEn
XEqCliPoMjPdkp3mzD2LwmH5asJttQV0RuiCVDxgzywMz8gEAw7+iA0cDOpfuXONRk8hIJ2c8ptg
bvVKEhD3EXjVYLloVPVBaVO7yf7kph2sFkFsYkS9eQfDbhCR0SU1C6KTHmJziKvkiGD3LxYWMFSH
KRHBXQ1ZuxBZwmpRaDivm7IY8oRZQwz/jHQycUH8Hw5zUL0gGwWG1a8CRFA+j5jNsLjgQy7GIscE
6ACf7lxoOAnjptibxtWZXwfUWtCC6vwzl5G6bOUgHCqk3PqOb2EWh2Vz4kZyGeXuuIXLFK3YweNF
Nzwxt7a1ZP8nbvVpHf58NSfYYFnGBZH7ByXJ/3E809zU+BTdsF8/lBDXD9Wl1Tdb3ROdOsgpJBGn
AIEgqWvQt/MFg1IiybYmsdKPn4YXLCSRkF9Zlz97snG9tIh7VUQIjWbi9eHZKInJcoqG2yWtp+91
6CCfxCuOUVgpW/r8W0DkgP+aPX96K60q5B/ArUgCCEg/pWaGifueXZda3lHHWuSkTDNyyBziDqj7
MJQJzIGdEVVgHDHovZk035asohNBeSEr6s6LMVgbw0uH92VA6r/zrRhpWo5vrmsGPEVul+nsh7NO
UNKIDU2NTyI/6jDhkKQ5J3ZObCkkf4zHdv1sqgH9hMleVtffapNl7/ir5N0OFiGY+By0c9LETpbv
xWKPzWai7HmY1RtQeutzp5xcVBd2ZzSYGKBcWI8P7MWlmo1LJWiH3RvbfQU6iV3mZIVlGy/rjRn2
IZzU0f3qrJUKV5Qs4ZAJqgHCaV/k8TV+9qYyoblGjq7TbLV+xgAQrY0BFHMQwtxqc5fOhqHZkmnp
WYOwE9Rh9V85K1WxZP+7YA9f3ow/uNUlELz0nFVu5m8SrmTWXLNcmYIwC2XqeQrtez1ifmicmfTB
ki/+2p0e/2t1FWmF/Dt22ggsjqjrLr6FRp9D3EZeGc/L5NVaKKfaIJVb4q7ePEfnpDd1DuTKm2+1
osmFN5j6dhnP9wYaiqYl2CelTJvd61KiP7alvyXO+PJhT4N5VphfJhS/iXGKNWMiz/mSRcqZETqh
puXeJMQfgG64Qi/HJ1sUEAl70Ry7nJ5X7MT8gWyqUO/Fnj7D0YPEvw2hUiUqh7AUahda8Se2Czn5
idHK2KkjRZbZlicd1jTW0bu686mwRMqET3cIMmMB7zORTKK6shnQQRAV82Qv80Fb0KWeBsuX8Sjo
Y6r/3rA2Gsykc2y61MQClnsRBLrz5qUR263ldJJWEM2b49Q7Sl338nuh8ynynqxco1qP0dJyxfW3
hvDOl2rZrr2ES/umQRS430/DQ6v5rPbGYdco3qK/ps/Q06Pt2edjBQIHbO+fx7jwZwTgQUKR/mHe
HwL0zYo14TR/WtTXi37TBtAdFUm/lSg5asounmNZ7gjBgMgXuYRtM1T6JER6YHNdzqiCJKT0ixGR
gRiUTiSSEWWDdmHOvNKe+nCI0ooJBtXZe3Ydsi+TyJOVjSuYTvi2CSvacZwrg0fUMLflX+jmCunW
jSISZ+yFreq84bxZ9oP4FC8LdbPA3kE+iNd1fcDLEVr+ywFLK8kOAKLYD7XkkPZLej65Fw73o5Z/
CVLte56bRoFn888hcJFej2imTOtrcjoygEBZKJobY6npFknbHnsCxcBExES1orgeqL/SiNuHTozc
Y5ZDeI1feCJYCnF2ipd7ucjxwDM+O73iReA8tyliIB4H/J0l5nBPsgJaH+t1Uud4ACQWm7r/ePBC
CSc4dCzD6JYIGbWYjs0xF75YPPZ4ffnHgE8rTlWCv6bonvz4WgA1S+w2gNlOeVrfzwahgP0lAhbD
TNGS6/pgv8HcTYb5GOCB85QpCwyHKHyCRjd79jDBnQFMpv6JX8jCyc/FSlzP9xzElvMQ2RKZVxlL
icPpxRWGNj5PqZbzBSC6O/kLbpeS9JzojbQn0bDe74I/9lFRMQbj2z7yw0ZgctSp8pTBtCqUArCh
yXzjxv//f2RpUytM0yQFxetZkmKkAFldlLFwThdVNUT1bnzkNOXQSeGh4Bh0zNqMFbCS+ejZu+3G
hswm0dMlDQSup9DSkcbhrwcu8TtAKbRzIPn+g9wBQhJJXBYMP0oWWACZo2mgaVUMnkzUsuAGvkJa
wxqEPKW225fTRHJpX2Ypcu6HbccAOEx+0s9bWZ/cagVWdUTJs+hgzyxobAm0NZM52kVs/nm0r6aI
DLFH2w63b9cttKUEh3TuEgyzqEwfwPoFCuQpoKd2sN6CjYczLbWc5Y69XsJSTw7k955YMdOD00QZ
ZyH54EXlo/N1eT/0GRhWKU8jzBcd66284E8pxsW3630yNeRApHNh1lHOc4GOcmniAgLXIx8oJ3Kd
henKqLb41yOsEUnNpYTrn+HkhgJbUJbwIHqnsx/mqfgH18GsM9QOHM6TsvwBjbqsY+JoDqIBC6pD
xhdsZX6wk1EZ6ViJzAVZG5oRtca1qrH70CO/LwzcO5CnoDiVe5VTpiYADIPosBuaNYFg5CdGzFNn
tF79cmdIIbtIiUQmgoaY01lu4NaujmiqPvBdT3SsziX6/K3rJ20fn7/PCcGkiCgQha3s48PdM5Fx
myA/6avli59D8FQF7AhQf+asJmsZt1qKq2scNXj3iYg8jAcUjyL6vjYY5T22/B9mkcOmGmkrQx1a
GARiihOaQAmX+pO97ddPsrFlboYq8m46HuTXz8RZ//HD2lZ14pqpez8UuySs+bLItoE4Sg4S76ei
/ni1KeRLerlomxpwwfYHfvvXxF7ZS6hW8LEZHj7AgebwAGc/LGVTnn4qRMhtYj7Cg9NwqNWPOfE3
N+ealh2TF19+EbWp6okdgt24u9QQChRfh0lSFhca0VBljrO1vQocmTDQkGzuP3XsIuVLil6WgF5G
5+uzAZhuPtEXBXZzkXQJbccx3i0RruernW04el8BEbTkiFfg/jW6ttopYIwWYWj9tLscLD7sJPI+
YT8bRPGVW9t5nosJPeKcJz//POzA2RlDPjEIYI9cf8ciGVczTOKZNtAYAx7Vrs0SGLnypKMwEA0u
zzjGjtwPTMhyaHRMPCSO7yxvl+vpznn4sLeLzy1N5pzsNxy6k5L+S9s05SAMWuPb9B/3wYiRyJcj
XHIqCuHLXm9gMKQfiTh6tEtUFNZlIeY2j6oeaCKMLNysQBTuzodureF6Eb86mH8yxSUvCfXJm4b3
vKMHhZqy7ipYNbhN3BkZ6fXj0G+J8YY+TDxNAkYxU5FSfyYGBDa+dVQFuhpCqOvbzPu27RP4lRkQ
itvVrKTjZwKlDvgdARrZkmlttj14gQo00xSYbsUW6HC818RvCABSxUETLmWhLxLCJ1Mg6pt/CRSB
EuxrG3xP/IAUHX7aGSKkXWNY/WwLcXCmy1byZheuSYEVJg1qfEtD5jJlv2FoMyp1G5btdxikn6H0
oqRrGdvcNArC1LtLzBVB4YSIM6X0pb3er6FCsLTOCGm5G10NUXjyv/7kjbH43M2zRsXqGDHURRnF
hMeXluu8Fd4fdHC8o+k0MjtrA/qDIy5Es1dXPsjVKwgW2kjb9N+lbpXe3EHuLwPuLyNJUudWUrh9
ifmM15ZHYN3BpAQqO/VurRfziQgpod/uQVo8L4xNZZ+feyzZ6TodqWVngDqTciwHaC6wLwOsWbA1
FQS9nUsFmUy/9rsoCIuqFzAW5/lXpM1azTrI4X8E4Q/WAlWzPMarQad31aRH09zDsttOf4v5IMa+
Ty3yrynCg8+ndLQ5iZNRQjwTRv05028OTWuy05IUZKc83QZWN+UmXyRkJqVgBayJX9qGAq/PotXC
ucN9QOjsyTYalG1Es1Tr+gfJC1+CMN1GU9Rjlits2a5nW2qSB0JgMO0W2rTtnjrEch4IYCC2UvLF
qqep90YRCuVbhFE8aPwYT8GMIrAT7QDaeQ5OPkClAxhWkt9jbFKXySL2ue4p09gV1+8W7wePlvbO
8fiYsM624t546oFnO+Nga86qw4f4lK0NIPK4ADWqJizvqcLSTtIoYRrvV3F+uJ6ozRZXvSrm7Ea2
IHtDtabUTIKQk3JHPeI6w6mtbGeo1ICRLoqrPobVHUQcgeZwETslAy3bEw03zTqblsvw2F3BQnXG
z4FAFEtfQG3hKRfUsQwrQzBPVlmSx2M4k5ICr1wN9eoKPzfdRZjtIwAz2m4fDFBnBsTj0d2uucxt
n+tocSLXA3fFkAlkQ6sQVX0pEMefLRTvc2FtD2tQLsz+H6dF5Eqzb3H0uR+uuuthOU6prtG34jxd
HfzxhGSt/b3O0I2ZoPMJVfw+OrUhSkO4crXGnDffxytTfiN7mSOm7mHiNTtU9eoSocqH9vXpDfSD
4/j7uG9J4toMr3btBYF4ZBICL+KVXmG9C1x6uiw7K+45wYGerCLwRypsdmTeTJyQVqyi7is0VYXw
GWSUbuEmaVZXyZKRLm67P9gjKO4b6aJvlULOMeY52SEiyNEhbmOOWoZgt2iqJGTAcX2otIG2JW3R
pIHv0IXJmoJd+RsBjXyyd2nk66nWPrF+h0QLLWz3p4+pJeYnTLpFK5/UtT34QJXdwYwhH0vDfZb9
l3gi4MuFSIUmHLdnOBXMtdOkXAXzuLCaZKWaYVcErxcPlMaSoo468ewVUQt5BJCDoLQhnDd8+upE
4hqs0SHJ3LYj0V7sbXY2eZgNnG3r1nvp88z0vn99eIpavK5bSZBqR+C7CIcrpoEwGUcNfyvMo3mq
XsAi4mIZya4N10JLEag/1MJ7ZG2Lo/cInAXg/upvV932cCEEI5x7K6hmYl/SA+jhs8K2Z5uD5dYG
FWT6lsIlmTS2uLW49qiVbKupabEhd8aF25/VysSozXrqIqC83Kp7uv601wqnOlPBqSOyIUxied/e
RbBNOyn+SJHDFlPD0ijq+TBCrLZEepEpQXyqnd5uelYtD6/0JYakpffMZEx+dIaALlqyKNWJkQ7c
CiCbuJVV5CQUEzG8/ZA1VYK9PrVlHj01LEf/QER5DWbvwmpGnfMc2WYQU6+xuuUmyAS+uiC0bh4u
yfo1fBBg+weGkfGXOteodeT9G5CzczgXlqAr7BCYiwJWTIGAaBaruNpNJIlDCbGEUpQY9RLGGxII
jx56as9UYWKOUwIYeUjBhDSwRNhK//5qfGUEZsuW2fFyIPOIqgVpkXdGY6stlECy6GXa5NwhdXPQ
8OSDpuXHfhvrLrVEoKCai1L1LHmtDSDJTLO4MPFEaKjzopgDwbTpMmNgjdujiLauSSiEDsdKkkvA
z/LE1P7oJFsqvhDPxWyyJ2l3vpiLwLJ6fHC268kt2LqF6FI7db6rTccPg7UX22IBJAcMu6dyz6Ex
5q3E2E7bvEHSoqZScfF7uuta1RVqxfekIVXdhEYGIvSbsgog4aIFx89yuOQz8HfmkUO/nHCgGHoD
+d0Dwy0wcuFIrKy79YkhLdHGcwCg3UcZmZmAJ3/H3nZQEvGFlB5M8uoI2ZNv9PDcFGS8X/UpMC28
3lQb7XKBN/nrCLeuHhY6pX8iTo3qcUEP2zEVBN4XRIO/dVHYyLbAzeyIJqVmKFDJFI1t9mEN7Kp2
x3CPmKHqtyJkat+Ph70A4haRGVTWt/X2L47qWvdLRwMciQ+2Zj+ylsuIrIZy9rOL13AtNtRy2whl
M9UvweUBgZCJRqOFRTRTO4vD2XrMqzAQ/IRuyrK/lXrXtpe2L+tZrqTlcNMBttz6LFQ07r8Ktson
p9JTYyZyLEkVBA8QQ6WbKfXprbWrcJs2sf6QSnJTvyHzbbxZeXvG6tRXACiwe++9gafDehSad1qv
Bfm5/KuqfVBhs/adB8BMiUa47ycTLQvtH6KNx1Dfx0d0n2aBt25xCLFaIHkMFr51gnZl5J0aw9mm
g9YVY9CZVbu5kcn0qZEKakjpVBapUGuo2trxzOhZWvcNQXzSk8PdQSRLycu0H/HyV+qnkgRq9U1G
hMjbgaWd3sGnnUyvpavmVp8zuEoGOdosCSXx7KiueuSNaTW7aW68UqP7CPV/HrDSsU0DkqFTV8V7
pgO5+n/RjxqCi3Urpo9vFbrBhZvoYS3MGbRbisjCbA4cipf8NlA935HYOq56yAsNNjKsAHhpAKMr
Uh77sJ07RSRb/eL9PTmG9QelWGFURu8ahOvBDTUghqj3O8wGVD3GSwCOlcxHjZ5fVSJpaS5cE7hZ
Om32Yad8TLLM5Zd9sAIgPJx52vNTfWWvARiFRriASh9kgf6ZtSsE+oCG71HGRj9xsKe59BLGpJ+/
LV0MUmfJq+UHn9VlSgipJpMYKHRnhwtio637t3DkUSP+yqtaox2wVXPNfH1xtnQMLZ4NHifZITQz
6lgTRBTSmtxbwQXO+QAwUPwP8OX7OJJTzVcWvnoFdJD8zl0I4n19nHTFRL1F1w23Orm73/RHLOvX
UAzO53cs1uZFltE0gB5XEtFIn35tcrgKvQUBulrdotS7ulwdhWToIGYt2+r+vPU/BJZcbVQMCS8q
QqM5Dh+3Zp0VkhQPAUBynAHga14SsqFdUm25GqkH+i8SZuOTPf+F6No1d2mDg94ZZoTgAjiyXNQ9
SFuATx4YdKSO0Pl5ezXgRDEUk9CfDsfttdHzTYigZ3/bDDvfjvBUiptQ0wZ4OgqZJLi0nDR6nGGX
x63keIeD2EjAg+u75dLqyvAenhWUox1Wr6ING22IG4SV7MnEHb8SRw8SGnGHe31iltZ7LS4mvtkV
BlY3R3JCna4mJFu52StPmy0omU0aWcK6189HAAfFYEDPLdE7xa5+nuZge0QUvOtkr2gvm2jbl9IK
oLwI//w2ihl8YFYP6AdqnqGiw5N6nAM/ov2+V3nhv4+zD/r/LLusQre1eCxIddbjxvLYJVy7Uf2K
sjmsRZEZH3DmxIMJmQU7UEwREzx6Ts3FHBDB/mDCAx3Qsh/2DcbujURVRyw3WdQfOXNXN41DaHb+
/58ZW4CjvuUOx/WzJirW4imNdCGcRag+3+oi/TO+CAH/dkaOygGLJK021pFE/srpl7MOXYuk+eW5
gkcNCRZJl7nyuZ231ws83YLMY769XDv5GV/HEz+XHXweVPSJTtgap++kcX717TlfMOwOfG18Z7IE
FgFR+H0x3Cck0iaY51IKL0vSMgEYElSoE881iTI+LQks8iE9J49OWgF/kf1N3fmnAk4SA84/mclw
237uCVrzmbSXM+8OPBe2PauTeUiQHbkh7gaYuKuCtYdp1BSkqD4lsgMyNQK+s2dzhY8ubWbxG5v8
ikpLpSMTd/5ZjYHzeCIM5fSXYYh+x2p9eMafp7VbtEb+lPGQSTZxg3Xla/TfuSmdSizTsEwLzMd4
Yq98a7O6yOmyXBOE8GsS+s3Z4jAmrnLM9589KcQ22mkpAjMTCTlXkk7BctmDMyz+AlIg8yttISEc
n+zDPHkysKMqDs0ETIcokkuC2NnwxsH7fLFyjoXw49WnTdJxfrp2fQitvm2ift8b+EClnop0DMX0
b8stMW1nQtVdx9JZlADL0QbCsUggy8xgub+ZvWFyOoMH1jkUt6q/VjfhQyJCEkSClFe8Tz1ejr8x
epljKwYo2EuQeGmeKQZF4lTRB0o5jbh+59GZjDgaesuYdQrfkEv6GKFhirpfglRNXvvA1yTVbb4l
L4ogkgyJgptZxFHsK09WTbi/xA7KPa9M3uylIIG++dHRmBdj/BGp3cb9fnY0ATo9K2VulEcpJ4yy
kxYbdFJry8l70AfxxnaDxLCxnSowbUroSPR6jAjBqjgOsqZ3kmlY3JY1k5V6gidzqh7br8GsNCcz
b1sBEorQ/jLY/7VE50MT+Xvaoc1USGSn4DycTg8xfclcZQIp9Ly9gaMUIef/A5xSAFPt1MhlNhjv
LqvR7MwQkDc3uVCNa3uQIGg9Q0fj+/d7dbcfz0ObszfovhUGzFQ3BE5Cb9vKpZpGylssaWTIhWva
rSA6nTHtYGfe8NKKeo174Lk4HFA9w6pVrizL0yS4AXmO1q1wkRksFapUgK0yMcrifACZHY80rvUC
HgCnCY9ldIFUYE3l3AtzPEsuOXRJfiWd4+fviyGMJEnqX9gk4Ev73C24dKG2i4CIHEQo+wTp+M/J
/TIydIOnfrH75RI62r+GNCMO9Kcw9S2OWefksA1L+6QJolufBzn3P7y6iJCqTk7kSG78PjH5o6pD
RQw2ykTkVDmfvMXGtr4wSh9HLxIGhtdtxc8zahLrwp6FbbBLfeKIU2GB2MrGwuiVQkUoTuTwZ0ou
lVrfyWiqobJrdynBh4YZwWJOUzLeesM7A4HmGvs49CK+tBIh9RCjw8Q3RYahOH9MNVNBb848hzhG
Hrk/aeNj3RJuvP8Q6zAkAZK3bNJczwhsYgFCnmqwuEtSZHz9krUhjwvKZtR9DIA1/vE+cnW/hwGL
rFtyOUfbk3Pfso/2TsWRoX9QVrO/69FvAPBYLD49oDBODOjLozqw08SYmNu3VJvJ+nUHhrPvAP2G
V3OhJmxO8zjjH3WS0tx0tytw2zVPKf8BkGp0E40jry9xzN501k0p8hhrNxmUxajXvY977KJ5pTBW
3jzJuvsnndcfLZXhmJZcTb7okBuUBDf6rlQ7caokgqYjJZnauQ5m9++RJxjdiy6Jv3HfNnMWpOu8
NvoPWje8130W9CXyxkuD6FdVbEpUCUnXvR1qaj18k6v7DhBcBc4bINB3n5TolR2cC2kV1NuPqGFG
Nwr2l018TETv1TOFZ/KW2udxg9hoC+HWKKXzzxweIK4giCTuXHyB18b+AFc/40AIDseGwP8KIWkd
mjerndt7fVhhk4UPtYOu4v+zDxBxbUJ4XO8VY0zXljV85xgEKvS/O1NzfRp8byLyNuIGX106UOUo
EtlZXTSZF65O/SYbjpFgFtRkYGBUC65v1PepR49u7XoppPxPCelHF7SPMZYMuAlkwlL9rJ1GKb4S
K+DGlYil68gO8WLYetjTrYZw+ZDaMUb+rC1P9SQhDXllYjZaLZKzdhiOIGOy9pWPa3GjQXItnC5K
4PQLjc3vxRvej/MawH4xFAag9PMAcKE3/Xh5fFbQnV9VmRiZCFwKqy0UuJxUENTk1n9FnhEiDBbj
uEHHZ4YNuB4FNs6TcdSp76EpFQ0FJZfk037HjAE5UQPUjpYkCjwouz4yMkx2msTKWtBFsi+F0iFk
2aO2ptcYD4YRaRyGG3p7qCmyZ443XLdBc9Ga1AZLFkMJhQmrTvzpqeKR3+u8yn+C3DLX0h6g4pzl
Fu16A6w+G+rKgNumPBKtFQrXkC36P4BYksd5U2UcN0Zro5uCShGdDiD4R74z8UtbUPAUKkWYnqR+
bnRpSiXD1QCa3a3hlXSQ4ft38RNGFseMow30r054kyheh0wkNC0WJOBmw1XPvjhOJdjh+duA9yYo
hS0H3zxqeBrioe0gZYiImhNw4PyaIF/xCQds7NPlgcaLVi+NTxvP3bLOeK2urqWFOuqrIhX44kKC
uEACAalbH+ZmFwpO7T0HsKDk6vVve0s65ivnFgMp2PnjAslXgnZnPWHcI82nxOobq+0hRFe3Avv9
6NKGZyrUx3Qj2NoaRRWLpseE++JIm1D96H+GFbqn+Ms0xi9dbIdlWUgsmMJnU0xoXLPvbWCQIemY
djWtLHhGhrlPyBVur68wR4KkY5f5GXJ8FpLfhy1L4wjLOJ77DgoUYfCeZdc9YrTGI+ZbvchSI8lS
Bq8CDiz9pfivOKxK7aCFrqtqN35AmAjjA5AiZN8XoN671gqK4ldnQ6CLZ9KEPjUeXLSRtTZRfBYM
FAoXuDdcf4C/ZjnG0KqSWBD5E2VbfxOBErA/zroYjihwD5IzdXPD6yB2K751gANwHfFFqZs80XDy
+vXKxHVTtkGYown1VedyUmJI8HjdYYcp+R2TtylXIYq/81mxDkwNUJ8u9TBsN2+2ETL14LhHPmXu
1J2ZIfintR5I8oFSRpb/S7sTefq1pA0wC3f0jkWXsfepFZCQ6xLrvKHnqNccSi7AOwlkmyZsM2GA
L4/qiZUACilS96zFrd5ixIvF/tawA4VqUWKn/kvtFtrPTlatTraAeUYp3YRwPp8QKzq/MKxeYD0n
Y0n1hAedCM/AZ3LlWFTN+Ru9PcBPoxiQou6OeyOxzfPtC5ic47COjc3JbPDu1KSjPbmOwLSm+Mny
C+HKWpoJ5lIGohofTzaz4xBVoSXW0ywaAKJ3Hnv6BS8zKkSdv1/sGuqyAEXkSHvorMLDX1HZTTG/
7t2bvH5AZkU99isOCN+jMxjPRDbxH/9S31Z7UsFVei8zoa9xu0W8GZyJFtg3Ohst43of6oHlD/1p
4iAiNRlUFOUPg+vw6RXQN6f6guVqi0DAeovW9BxIIQwucyzwVgOEfq6VrIKqdWZ+0/sW/wBS6Ebp
+R2XixxfvFWU0KQZS8z3ccu9MxV/dTGegos2OWh6ChKZ+ozUybtyDupkAIH2aN37nC3So5ra7kqr
h5/tdt+4U+DXOdxh7AUSWKl65ixJx9IEvaH8LB4dB8U92nzQQw+eZCIR8aCBAo5NzGG+UBEpQ0oC
Ck7wnddCl7/+buIg0nOF+V96aXOw3GPcCu/esl7F0DWSu7zFKoNOMRsIPap/jC6K3hIq/DSD56+O
jsM/DzDCWOzF4wAtRCIfgnRm589JCIfD8vfVyr0zYb3YwxYmnH4WrCHToYn1k3aajtPGyLmz1j6B
LtVW+aovE23eIt9ND3vtDTcJ5IktknH2F4yxZRty0J6WVNsgwrde1aVDC9nG4bvvjHdXCzygHJm0
0tBaUWpAVSAUPcyw2mU/tFs4GHOdoXAnHjSO/xvJyx+zteOrFg+qF2C8ujQ6Kw8l+96SWmqLXF0/
s9cCK4Vj7FUJI1Vh2Xfo+qlWGgc9nHgTAsvAlBiS9I+n3c9bwtyRfq+aNyHZSzNZ6hN+XAxbsObz
q7u3XctguQJziTh3UUo4TjG6iYyfu95esPUX9a/73nGTjpHc7zi58fTWxwdgVTfNo8Fiv2VDAlWi
mt16Dwc062TkAC5mEWdS5L6xhZOZAUyF58YJMC/XCxleHLRLt8WTR1sb2/eLI0tw903E+lsmVHjF
d3a78663qorXMn2ky+7kHDx1WvPhmJFXEKgJ5h2zpPCeOcQ3nfa00cq3RXffikxE4ZI709eP6zz7
9vXngGDZT9BaBM108WbeQk+cpRkuv//hCzLNROojaNPBEEzgNAxUeR6LN9GYEUDjUoV4lowBkXdM
AnNaPeygvtUnbujWwU/HXh73+nz6m8ITSd6k10sE4aoP9Jq4HuaREVv3TK4wyHjIb9bdnH921Vdc
1gUdsj7i+8CybqiEIdhk4BfXrk0wniRbgNLzWEsdjypcBDCXh4k52KgodsXeETdVSqVfzvtHR6LO
1FwAXsSAk++cmXMsmOsGPt7qyRG85+WCPqOHZQnRnl4nmRqPzRaUnaOkLa8uY4vjEmF5zt544iQR
xzrl3Tc218btVEJIA4yfTgkXJ7wwRrSoceQ1SJsSONV/50ZJriV+t51yl4RzbqNlEJOlq21on/eC
/IUtFJR0/hzwxURF029Rh1rpEi2paZ3MkSmXgORgsPDLGQbnqeHkcgkZ0R6JnHxqYa3LAllQnT8X
qnbaawy7cTH2+3BmVn+yI8NG4v+lgf/+kZAsCrfoXQA7dwRHuzhz4m7hGWkA3DNz65L+1+63v1Uj
SWuPJ+roEgUalPDtpO43qmejh/gfZ1rzAFUBcGu3zW73tvoGCwXXimAywzBbOT74YXkHA/2uEWyv
GaBUhioCUxl1F+qS9o3CZHnMcgcZL/8VuNXi8d4hixu9o9ETUiUJsXaLrEGY0j9wXQDgXl83fCSZ
7DT8mx0fdmpsgYhx3IO8xmVsRKuhZs8mOOizv+0gLm5XKwB9LJpiIiF7urGMRHrrWz1qPz5hRZpJ
Z3G7H1d5/EBg7pQqTsUJb7hKfS45RVPe83Qr3ISpe0YNkuzMPxFp6kEpKCB43BGov1RWS7U0WGRi
0yg12IVwPa3yEkgkBs+el/kvUc5s3OELC53UyPkhe6c8iefz39lNUubrYZ9AcdOVdOzciXmzIT1W
THDVLFYJuGLYqPUeUXW/U1l33tE5p1am9xAyTRF/Gng/XQh5RpzT8Bp9yU6HDdCE7plXgEuzDgA8
h6E9ryWm7/KFJOJYGozmHmEStckJTtPX1kDqSdo0GWwWR6qXRKcurnCQa04dS/sW7CqnmC/qJ/fU
1Pal/llTQVT1QoJuH3TYC8Z0rorNnddANiN9D3tQsLxU9sG9w7edMAV0AY+fnzDH8wEmJCm1ob9H
NrR+4V1Hlcxd1XOVFQO+WzzR/xwD7G2C82lUx+t93if8tbKpP01t9Wig8QR9FIgw3LHka7Sm+MD/
X4Ews1bvGb+eusFsqjcWxSCKd+iP4fGslqWMqVKQXPNCA6+j+pteBS35Km/CU17ht+mMLhpqIVGM
PVyVsGNY6yiN+oMviHHoUJvanmVzhxmw2Qb2jGE937FC5V3qvarfHCYGMDwQZx6SxEfV/WQNdRm9
xZPLKwDWjyfuhLzoQtWMdUhShaTForpHcwYLLFYUpsaTetw02A+SKQzHQK/LHHIKSDKA2bvdxx5R
VpDssKbBPnDUyfTJex2KYHQVO/JLYoPvV3MetCaJ0ORnfFP+XRer5UoGT6Y9t3VeFtXfDbxrctcE
t/LEbF0V/KtiOTDgtfj/HCpTqf8ZmFPeJKTvzf5l1z+9My6w0in1fkd9yrqEmAdLF2VP+77m4rOU
YXlZ7NOkmVmiOQGepQ3FKPPF3XBlZzEyfM+eyzqY2aaThx9t4+XefbnSGJo0R21fJJOnFOBYjhbY
oL3cu9WJUE2y9OLauzpoOW8xPrznUoH00hjeROIF2Q0gofPjTmhyQH+Ae8VgywnDKnLdwmMp5SEo
1e+9fj659kE5yU0hsWfwz1Zko6Bd9a5yE+II/HXU8Fo5hshuqZUYM3C1c5psK4v0k6PyaIunkEDW
PXPd3MBDmUaT1XVFjskbh4AKSXzB2OqptikM4pDUJSDW9tuWk0RZ0c+5K7/DxdMxRLL8zJJod0Y/
Vw6gZRZmK/f8Ek2EeheE1gTe9q9KkmInoQH0vIak1aNQ/XLHfgb0Rpc70yJlxms2YO7H2TiwQbuk
PCruZREapeMEelN5e3OgalkAXa/1mq1ZAe+3UAm3L+ANEg/XgTA3WlPXDC3+VsARdR+d3+f40vVg
KTVwE+wdlDvCc42dYXLQA8vkvV2jtPqJ9h84qSuA/l3VB7b/QFVcq+MRY1FMbmCUCHpxuQufY1BX
8mmzQ1tIvHDAb4VTWczlSyblftrAxXDvUl1/PsmCb+KE8eYNNSsDdGy32JBmBqcr0RkE2Ve9kQj5
ytbxfT3HQGpsJpy1Yv0Pc8ypRHq7uvSl66NBdPI0doKZYdQF3swQNr8yDs7nuzbrsy7LLQLrsmoH
elNUc4q8S/4KvHr8+WAA+YAKMR6EIws4dhYuJea+8lXCVqwCV01dkIvNDPf6rCKv0HJ2NPzhSMqq
8uV3VHgkP0h9C+hoQOT1OKY5UC720KbrwyIjNNSvX4Mko5ZGhUbdM/mhq4TmQjcW4ej4g0rf/Cxr
9exXu408TJNeyQSvHo4JHNvLV9hFQKQhhOqNNsdizjTUhER1Duvnd1207lmHBbkHfKsOj9gQfcQv
egUkZ93d+/58043+iEYfmjchpz0h/cXhThHUOVMWyaxCh4oKVUqBcbUfOFe6OYpkPVT+QZRIbnzX
Q6T5lQH/vkZq1EyWPoYqdpre4GSF30NtzVSlGH2Xtmeahr6pLBnzchy7I8QNcFUyNJQfkCU6jiR3
t2pOJQsh1EEYjihF/D+yCd2VKKkLm/u8OZauLCzCoI+WwJpKEAz1S0KbZlsLq4cz2mC8n6qvY4CH
Wdwdbr0ohKmKTSR4BXgrdcPeZmSTt2EoOV1jdaj7m0Z5Q6QdP+mK8iPIhhxq5to0lvblybAYx8O2
X13OGeGtT/vrjNkUg4x127YUYwYb3Kcx182xE7pGcfCOaWM8cX+5X3lLf4BnDRRXPECEY2JYX5pr
wwe7VHv4bFdgl3hO3vK4jiVrC/YfFDvtnKSW/IcvqaGupdohDQGgPdFR4nSGfL1VH91iNWxlmj+T
7J55ZXnIk0h3WJMBlXRlOQLwRWh3lQZFwIDWS3DaPLUWYaqFCScNRKCD5sZi/5z7uAx08pLY2djX
df3GXYjWcIWJJR2lKYBQp5+wiN2veQy9OqxShHxxrkl4AuLwzUNJVOYLRsiyoo1KDSnxz+ear3ZC
TeBZv/xjGc3kFOKtx5958lqcYOKzwT6eRuTvEDfLi3j/kgWtvZ0W50NsbnfOAPLdabVjYHJaspKD
OCjvfSVPHEoD7uYsBMK8605yd6Norqj7OBky5ABc5tqM4zesD/ZZhHMjbIFKkj216ci1LTlcSORF
rteXalXTAyWkU5eJk3YOthBiA0DMF4xWaW7JednwPyFs5q7TK/ocu4J0vuKA/j14FNbIgjNb48PQ
Hajp/ailNy09PGqt3YkOibrp3E9fBe7Dh/hyHjWNzA4VImtmln/fxSccQKbIV0ItUKpJcUkIvOes
t1O2hpKUldD6oi+2uhhS3J0hq2+1tnmVqzEVI2BpZAZerrGrbyqX6njmcinIP8zRFcmCUG3LijrN
yjVvi3QikKCgXuf3GE2VW4NtTuOjpmaqLNI6xKAlcnWQ392lHDKFHUCAsGC2JBQNxPyaW8DyQXuK
WQIHqBr8DJXATiqhbkntHcAF7bcaeQiInyakdVeFt5e7Wi5pCmrjrhJ9mUjEKVhdRD/LrTqbUQHW
ooOmaj+sXmX1zXL2UAp5TNNtPVHd0kyAoCMqPXHwmQ0aVFEbFaXuwnMbqaOsEjYw/FQHsuY2tFBJ
lVT1IWik3gukksSsJoCW8Amsl3aa4zMAF+1nMvMb47aOM3bfonI0HVu+ofinuJ7GAiAUkJeSRhRt
o4Xp4NA9OjiUA4caX4BlTmZjygDroLStku/sUfjMgvD6XYtT2pFwT1MgRhM8cUhbYglJLCFRNfvt
L9s6FgiIQo3nbZbwiQ3p1T3bhacOMM3a1bUeCjIVP5x4BwqxxIaLzSqSYQiZcFZ0Svyj51K6qbfL
9RGk1Da1ygtfN3tSQkDxWlnT+QniZ+2mNqIdS768vIDILmvNJGptxF4Zd5Wvws4MDTGLs03ZxiUL
CBV7kqJ/AZPugW3aKs8W4z4iwOs+YRVUSjD9pLN1Y7Jbm6pK7BFQiOBp0ouNyxSOjfGK6ypC1tM4
0BxBnqa4jd4BhvEFXtGXR0/UmXNeRKNEUkUxcMWgunGtjKPlhEp2ctP2nLyuuXma7iZ3F00pcnrs
t8Iqffo6wZhBNmAqsnWTNhIWx9CAZZo8dq6hhKE5XhUs5HSac+g6hQ8l3p6XO7RqIyTcaumDHWBY
ECGjHtURdHVgJOjo8xDJ3UA0LQiD87CjiGOI7fB4XLGWRm5WebxTy42qT9pTZZz2r9liMTWbkc83
M3YUgHbGRXIM8B5mynC6cl0zUxJjWA0EbwcmJN/GSqNzov5VI9goTGLUuUmDQ1qXpiujUwcK5syk
Z+cmhkan/KxQOy8yUFB02+6G0OYEOUyU1EWxuOkMANHM4XQCt3wq8y3Bw9GKSr4bq04BrhW9Z61I
tiG17U7cnACc7hOX8fWKYwOtHjp9Dn1zuYdNJqtMtMgjbrzTD9I9VT1jUMhct4hRtd1f2UOJkgx4
oKmN8GIfEeoNmiU6Bqu83lh6C6O/4Hm6D0PAJlnLQBEh25YRlL671IgXWF2q10zN/eku+kUJkvtE
cUd+ry9Sdr1i9yl4fRxLS9rP2RogmrwOMnjzQFJqu4sNNnhukX0Vdh7mgHc4t3Ib1flPsyRkL3eY
aT7FPyWaNDT6hWXLfsB56ctr+s2xpGvGCfG8UTntuWknKPXiy0NfIVvmhBP2Ln4/Cqtfqzau0wFk
TtqBWg7xZMgx68qKefyabWg+KLLli/rvCdgxJuekfY81z5jky4J5CW5mSyrSTCKAcT+NJZD7z8Dv
hm3O+eturd3NbaC8sjBU7s+23Df5q1SW2xy83qf+vozRJrnfchyrlz1ozCpBs9PFR/Jwkd1KICZP
1Vr7d8GygeOV7BJU1EZUCY5TNCur9Hq5WGSmQuK27OQtP+h5O3oemBlbArOXgaB6ZIjcS6+YMjNE
eVhUm+3I/gOQa4H1cuVIUCigZpZBDOcyN1vEFf1pnOrVQZmCIEAg/d+pbXtNbU9LW3io/qphS84M
dlPB2c4Td5AGE0S/iW8cIv96aKjyvKrcndvJMId3RDcvSaOeR5F14vNWAGhVs2K9QoWpNvv/WNNM
e+XUNAykG1z3MjAuy/Iku3IzFZ/3LPBQitJIW8670Xz/Uu1fOzM71QFBQbw7xZa+9vgqkKsmXfMS
28xldtvGcXngkFVt+fuYSfj8jrOvcDFuN2op3Gwi8dAeF5FU1Q/wIbrT0TAeSvYN3keNWKr1bYSQ
GGrWUslUlt/Cz/iywBMaPjuaGLWwlfs0NHXR0+qw8olPE7L8hNfrKlrVk45jEy/9A2qv1CV5YbGu
K5icDGyGByhITYfHavIP7u44JGWla64nLaiXBmPTVx2ziq8dedAFoMYMkLDxTTHd6bj7eWtDOZpY
UVoLtdq53And8MSvVeGLedn871OK5t4WrsYlkmowYBYHV1BuuTe2omYz4yPYyEDpy3JuWFRkVYw6
GMaTabs5q0ry3tSXJxohcNIn1jCPBA82pReAn8Q0keRE252rD+f8X0snOR5FDK4+7lb9899MHLIS
6mXmUyk+NotCSSVBrC2SUSLZJKvnx2K3DDFEuJrZRAmBjLrVTL3M0BoSI/ejE1Lorak+eXr3zwJW
ZcZUseayBB0kTjrHF3v7Vy7BaFvY9lsxfgnkWt1duMMuI3u5aepGS+c+aNHml1Z/SUvzE9CS4wnq
xUt+wEX9oannNQ9vRZWl5pouErkIjKy1IeUWbzaVk1AHYBXgwEmmsYMbaRDOm1FVV4fbN/ClvvBr
BAOkM/UyQyRjm4cOXqGEuzCeyNdl2byBZc86U6OEAiPbfme8vCngcnASmNu7m5QU7N3Q4oo4Ai43
oPQuSX70WbADAgyfGgIolZ/6pKRnQWJoz0kbMz78HG5Q772VBtUVLeLxwz+wYPJvWPbh/OT2kzEy
2C2K+R6NgtLX5zABAHbYjFqJPv3jbwUOG+id1MeeavOK7dosR5Cz3Bcue4e0K5st31GADiAYPYq7
h0ruQeM56pdW1IsbUfDj3Uf3KoKdhwoQJSYfOxVvpWJn8coBKMQnbBTgcaA3WIe5zb9X1vi2Cogj
bePmHpHU8deG+7NdqTIZfUI6jFKuEyh41rYpvXcE7FWsaifIoCn5X+dw60BdhZqRIW8RR9PxXEQY
mXAKvLHTh7N0EJe4G8XG6m8sUyyLF+ei5MoSSgOJhI1SCEtXVnBoyfCyNhwJxSc8ZQrAz9lureK0
7aJIcSRih45lghQn2zBlUz5zTyalfY7kYjHnXrhmWwwpTVzv9HQ1fGZOTTIIjxerjelCsQD72VMO
ciSCdiYk5ZbHCvKkpe1fxaN6ub9L7HmE7d8cdKcaVejREu2N2lMwjDLYOe7vlTKfiJc91jdIuDJT
Z3t1QZnZ5oPXijIaVGwvJoqfRZrBy2nQSujcEkV/JpyECqbcl8CTtjK/HVVfso+SC6sPaZSWsQDn
UjuKCoXfGXtGIdExIdCzNc5FyzEx73NVEYX7cSk6s/POaBxFmuLDSpg6GGSvhG/wISxw4+hKUj3E
9rnNBhv/TTvGty3WfZwiB72HcPG/p3kWaigyuJMd1yXboGzR9bwGIrofYec54ubfC97wAQ+acUIG
xBghSh2aIQNdlNQ1t6T2mojT0EJOmyZyr452aSXF8DLfEArkUKZTxAqx/BZj49/3FQb71n5qdYIH
+Gecjbd8r4j/VC0r/AHw/JnQyIk1w95LcqzuSh9cspQiDRFHmA4qlZF7EjyZXANSh3pnVAsItLhy
68y4y4SpT4J0mi+BMALfddCNn2m1SHCXfijO9Z2tg9Qb3sz7pLsmcxLDy8Qi5sRXLgFDtQOVZ7aP
SdncHdwuJwgHMkJnurZOTL+itoYHoP485PVSG+fDLvzbiGIZH5HtnH9tW47QJzhP8wmB9RGcPa48
yI+Fny9QPmR+pnw0XqM49KNzaezn97qcAMsEI9IIpFG4KVwULkFZN2vs9dp5P26btp+xAeAtFkfs
byckkMqC4ZqkqVelp3McQxZl8C7E4xzgsutpXOfkYTK3m0k4Lw40Ob4fdaDS2Xx98U3oFmsH9e3p
TsEWuDqwz5H0khtPjTqiod2u6I5lqLV/IRgshe6vzRDV+p7ePHCMTnr6O246FZc+KjZ9EBu85MD2
qDG3vvvTxZxTwAAc/OXQsBEXyOZCAvpiEf/zmGbJHEe/k8gZEC8+6moqUotRXrdQaJYgBHpQbUod
GuAOmAe4v2vwbBNC92UlnFUsR32QHk1Fyv0gjpHwZF5m5t05dliKKY/hgP8hlBCBA5H1hhF/zGVP
wvAbhFYP0LPaglhfSv3Rgs+c9CqgVOwNVUGzseyLPVqPHSTxjWpxA1vEnLSs1ZuFvoFe0pwy+NRb
kpGOT1ez4nX6qFd+/vQzAm73pG5jyn45z7Mc6wqH1zsX2MOhdJpl7upqafws3plTfzNSBDfNiKu3
zTx0mVvb4fRhqvPK6NgaEuBfjWMgpf35bbt31rKVUpWx8TptPCaoF5rfdb7Qsgm16fdqoa3JVF5X
4HIswADJf4GgJ6R5N36OjkucT37Q1Z9bdzxVHUDjJ7VD/0j50WSMjf1oxMF88SYtI4qzBy/8xYP3
gJ0TCBPndRfyi33wk+Gl7AhGJMi5CR/di+1CojrSZGX2PLlUWqSRSlqFWTwZjgjZ74uWXvcCpTHf
nChZJsx1kMqqOuydsgqkJw5l+DEDyGv7oHDcwcZj6knsin3erf1dMDaUSq0VVEwHB26Lp5P/tTCa
gy1+0yR5UYhvRKkChnhVyDLMsjQAi//dakN7HQq72U+5+hQwYwL+aeObOjo2X8NGuFp/szfwp7YY
9epdjxSEK1rjVICZhsNz2RcsDE5ESa2Gb8KOAtvVwombRvJBk3hnMHZEHXIhqEYwyFFiFfGQRCGR
xDCFyajEuf6IQ+ZALnN0Rf47Egitp1OmUmmMyACaLxLauCjjC3JAGjhlmrb38yUC1MEYKs75sihm
RFN+zJr0FCaeTi71eWtwQQAJNldhmqblSLwL81dXqrbJokR4I12TzAwi23t2rNl46LhAni4CvmiS
DsE12Ml/lx+1aQzLEQTGyfLwmQQJKL+ZZvSwLmAZMExoQjGf1ahSuMJy+HTobbfDAnq0u9GzCAcj
K/6IVkHO4ybEUKyaVg3NjkqC0lBSvsypoRSfhIW7rVhr0q806qBpLnLBRtZwrm3Uje6CLR5p9XMW
13BuDUhSIKQMWZxr/V0bdmqEDABzgoX7FZCItqSj3lGhRPRqPc9akk5Bsv6Z5coKua0gHa29bHPz
0jgFYiYSS0a81pgW7zujGqaPZuRVu5NVgGS38n26hd3feUZHKOzkPnnMoxPXSKf23MV+Vpn9OZlP
9j2RdvjdgPCI88yOlg6i0s+kGf9T6oJQfHBfe051nQxiTkGyRqRNMs9mPB5gAdqlin7JCwC5zJDG
oCp244K+IAjSouNVcXNAAApAArqYRjqvBpbsU+FsxwTxPTEMB/CPSDmGyOftbfunxNpWhg6xEVOU
2z5MNUryIhHVmkVqbA83CWm1jE7KDslw5Dpsck+IqNeNoPyjOP3pH37OkL80pSIYO24wsICtIFPL
ut65sBhz+JawXwWcUlZ7MOZR9cb80xCYtyErAPlFww8kPQSFe1j3T1kPvyDvnPTP1BvQOLHiTRd3
cHbk2sTbrJsIuWhWeIaaF0/Ip/gLcp156JPgYPT8sjnO7XdSHbkRV5J7v8upamz1DrsScM4iZcRc
qwvOYYgj6KpnHILXXRv75Av2zT/9g18bPY4WrZxiuqlGdua5VrGJ28nmlUBlDEA/diIJwb1a1ePh
j8LGitPL/xbc9KBwfqaITsltY6Egr/XQEn7tVjqtUIBVZCwMr2nnZh9p/FRf2DSncl7G1iUVICvJ
jum2ZS8UTcHyb3ec1p6SyrmGw8ST/tr3xNB0Lx7qCEo5jNR1HpQJh4aiXsVRhKZ24Xy4xwTbkGMZ
cCIPXzhmHmIQpZW2aFErhONn9vXgD8p/OEQyAYchy4cghphWiWu9inGZbEvRHNbwkj24eWT68mg1
oohUdAIBNjIABb4pleANuKJHUxWWcHNu6wFfNRxjJV9Ze0eLaZxLr9x1Czk2EweGE5/EFHcap2nk
swWBKBFmS/XW6PAplWpmTFHMmvM4d9xFMzmrVk+0AnVLcUQv39WOA9hf0AxciwxJ1WyWrHNmHMEI
KrM7/4SGCq6KF2GopONCSV3XWxyx2HNtFeLYrhhFRIBe3o+xUZVv+bKny5t/bW+ZVsIrRJynuhWZ
1CfQJ8UgA1u3L4uQ1iyJUuQ6s+pALnbnZlUkCc5wITV0ouBFdeIAgG9dkxtKLUFSpfW2mlrGDSod
ry/h08ldLQ7CJwD/JUs+I8Fix+bszy4nO+gLlLdEUCRQeJU0JW3QYiAnXw5If+XeunGnqUMcUj/8
1dxDRiqs5C0G1vDsNcGCoqtL+qxjiA189/G0EI6VmZuaa2r/pV4AoI4ZQvvRZX4zHLSg53VzsSHM
nmE6wIHQX04BEFMPZyS2/ygsYDi1+Zui3rwUooxh71D47CS7/TXxQSsQ8El0Fg4f55YJr3uFevNZ
10/lQ24NCuVkT7UmYkAXk0SmI8qwfMfaQEla7VECZVOZd7+AY/6Wp2g4YxIX54J4TsTDdVlihH1I
v/jtUXLyzElkQQF4EB2udewAJeyPyA/BC2jwL+iyzq22SQyhYHVyYzoeKSt6eY+XEyEkYFzzx0a7
RzbIdbRzqOLFPY52wMpwDoZswwUgdm2RhiT+d90n68kSVz87SqCwyRF24psTUgoJ4xshfGnjM2wW
nC2j4Av7OHD5rNh2LHJYXAxdbaXZSobVP59qBWT8C5oY2MdEQgcZwmtt/ZWPup2GZNNvemR2Lmkn
5dumSGkXmNYvjYAchUOuHx1NnU3hzLogj6ZNS1Lh8dhjqhKHWEo7YLnrszO8xZgLNYX6S48ACLyC
ckNn+FPNUuw5M0pG4inoJwB4bPi+Bcph6Dd3p8mf7rBfggBHyWpnXDsPldS1rZ0YIwWJjf8aBidO
OwRSsDgYEWiaqhxR1WS2eqBmkPbry1m/RwEhrMNp9JZypLZAUdzQhCZq2D8ZHMKOul6ag8lcHWSY
U5wx2ZfCF8fQnHZsSYikOw/k4CXeY6NiKUf4eXYiOLoV7EUBPRpEPuSfPxCftaAFbxWRjXnr5itY
Ee8+LCYxsXbcoVEUuWyW14XO83s+HXZoXyohWlnh2l3KGT7ZS07wemtt0irqiD5wIBr1ePAhlXVZ
q4X5BkuxCDsgP1wcm+l3yOnBgCnbLHcCCe1M0z8pnntepud8BssNgh21l47auJJs3qtrGAI0Jpud
JTp4p6tgHqOythBSNkBfIXOXdoQesXMrwMhWQSY4OMrqpMXPHPuzPlFSgO64AJlKgCL3pVAwOQBW
iiJyZu/XnFwY3BNssqqI6f7czMf1M5P33S0orPY3Y/diYNEkXnIJvnVWeo9fmXexQxRylxmMGnJF
caZi97/iGH+Y1BV0bCnQeGmsE5ONuCFvwJ0XnuURN/RyyG33lDAqTrpvDjgfQA+NUxk+xvlpPibk
poBDbyU5FOlRxQE8oMmaRCsFe9llhO102nGpns+vdOqmLJYA3UPzgMutLK+DwpEEMSHzHpRF/OZ/
OCPEd4Gn1b6ea92EN80E6bUweqYcpb/jhjiC6IrD+8FHkMaOO2I6xRkhyB/PwFlQ08wGRsD5phT1
+GWUx/fIIpgCzXt4eTW1Fr+fK7eGx8tchjuOjEC02nwpkEc9bKxIhLF8WoqOB6Ua7YdWZkdVRc+9
M33xD207MYpzVVYaSa4yfOt48Cq7lV6ZVoql/PErURbR4+eaDw2K+UxkjwEMqXsKDYBxzk49hgJ0
z/uNJOc0Kv81qWy3oeNBJ5gaId7nIPVkPXjQu9JpSeqgEgxEb6TDlncKM6HmVpR7K8GNA569tvyQ
oa+oXRv9hEGkQ1pQtXFJ+zjbZRb6K6AoNxYCuSAIgZap+9K4lbe7kHuneB5c0PSGEgAJ7UwK+hu/
dK98jz4LVFY7nyoFjpfNh1lWYBv37mkmSGp2acbdHGmrtb5o/w4grFN/lm8G047MCR7IHAiQbOi8
R0OdfSJhZ6ER557LXPGceKwdQJByMLEe0MUFMu27WTClLqFwa/PNZSlFxbyorOzQQIlIi/vr5PIG
EL8gNOGPKWU1JYFLcN2CrRg73o57cRW1NEr+YIaNZVvmRPCRAR0k+CdHk+AdyaRwEP3WrRdu+Qq1
ckGmEonGygUDaxrgnANaZJIBH7KZvr7tEHZsN5udXn/hKydgSuaFunyqjAiBC8QbsqZUKuU6khds
nm6dnla+6hXXMKyR737s0hslI/lxnpFVx6nD45C8b+pk0uAseSDXm0fr6kYer+/P5fBm9ENaY6uF
APwvllUSKY4suOFxC/FNMPoMnqnQoaumyIhy4mcMZ3LLm+gCSF6xhIX5bd62fjmp8vn4/4mKNlY1
SIJBJfaSBc/N4qB38lDb4RSY3DKDRCY2N8WZDpyJdFbdg4XBUrfQ853PFcCOK80LsRbScb0TSp2f
8cnmtBj9P/wCgGIQ/ciQPA+Su37EF4KXFOmpwBdR/ZKWyKPuIIxln7Yg4gBqc8gTMUEDf8jmEq1W
w79EcEYBGNd8fSjfPpRp85vH332bNZ/laAFAwzzGRE/SJUqaS9B7piwlzMbiKGn/JXYQEPSaEZTJ
ff+Sl7Rrd9BKJcslZARRJ5bNv45lO3GIeclLPtV+yGyFnsoGi2S0Kk9Uxpm2W2yIXc1NYPpfs/VO
ppxkljC7rj8d647gQ//THIgzQWT2nAsJ+BZ6AwKjP0BaumBgklDWyNTM9Dxz7Wk37cdT4JDCYky/
oKcmYj7ncJlmzSKD8DjvyHP+RpirEeG6p/fN0wn51dsnqCHIEE44VL69TNNe3SEWpgdET8w+Y39e
KFLXr3ZjyTcG6oC8IdaV+4nVBrySIR5BHEZuPrpybS4rzhCOW+Xy+/LMfsPy4V+hTC9lA829A46U
iDQk0zVSNuomi0e3HjP2N+eMK2KoylCuN8z95R5K5kMM0JeazDdDvpVK3XGcHKlu7LYw6AVtMHAE
Ve/UzDyPS1OFLwy5HibsyjaphDxNSp2KqKLgoRWIzG8/vXtgOuet2kvQZZuN/FmKLzNIxLR+vwan
k7IMSpoMzpjz9Mtr2P1F4vdljhoseLPyOyr5DIjvBr3Z7HWYg3GZ4auI7wZNoJkAY0OOzF4WNS0J
WdWLMfAtW4qZV9q7VpnSDadlqm1iNGOw7HgEb4u0FCZk9tQ8tinV89hQ7FBbKR0AapJ36Trdd14d
SNMmiD3IEInaUnlH+WYvaGPFdnJ/4h3qHIollpXNyBEUzUw6QlKqdz4rs0xUQFEt8SHbvKLWIRll
8cDs4y0tajYb7lE51oizLte/pRgxIHAuM+4X1h5K2Ir6ILG+QV5Snt2Qy76q6BsqfQxaC3RRPsPZ
k/WE78qrYvoVkC7kL88SM4n1nQWaPUWZG6OO6/XdMQDe0eZs24u+1QctpjFcG/i45vaDTUKrzpk/
3rawqlLHUt6z7Ae5Cy9Edp0wrOkylMYtNtEuY5kv8FZXsAiTcSjX5ONjZThGyD4ylz3vMby/YBHH
Gb08GXDusizc1DP9oK/tNHfm3gYHQNYmT1mY5NuCOSGZFxEEVUGZiXGhVhecmyEd/z90Xj1iztZs
nqsAhz1lLKnAe0pLij3HtNUXc3LWlC5yQWu2d2FfxrnCtTuBawVrtUEjsI+mv2Yv8GgtDFrbSjqO
H2Igj8eTsp8O/TOJq7zPtBXzjka8lkSyJb3ijePkGUM/1n7cIr60FVacY8byukBxTuSJPG1DrHjr
wlKvgOBjAqZ56WRlUGa0F524Jrw2x/7yvqfpsVSfrMNzYaeLfttmZnwksaQcjNwWMLrhZumt9Zj5
fttrNj+JFQHoh4tWRBnmZJrqr4UCqqvyDvR+4KJQhnFvnQy/ENq+HBAXVMIj0/n3EZiLwXnCr4vO
tJNbdqhz6R9tVmXwnljhikeR88Gz8z1W95C1Ud8u45PGUpCS6wm4wPvAxpZMKvNAguvlbKRPNQwW
t9PQUZ+9ZPgJk67p9zi9edeSwW0tKjOyMSKCNnI60OzFOtRI+mQsigOQqStsfBkMrC2FtzJFBPQz
wYBb3frbsiP1kYiofmkUNrRSVgVrevxAdr2spvzIMaBOlY7wtkQ1UUKC2Ldvf39Tc+7p53oFSumd
z+jCuvV/S2AxGkXzGlPlosvtwwYwKwEtC2ug5DL8CnbCZ732g3IB5WDf8WkvY7mQ8fUL/iqUCa7g
rNmY/1PeG13GJ/bsVNYecuOayvnGr3KkwwSZl2C0HSmernocbEYXGcq8CoMpYq7dJTFJ7EKX0pLG
nUMAwBYV3ZAh95Y0Zpky/tYdVAmbH4nwAUm2LR0yR3MpGC9L+DetIhNsFj52T3GOhJ2nsOgpC8/r
6Pg3Gqmhmd4vGXM5Y6SPTvoXduRNqp7sJHeiUhwTjqgy80HpaCqa6Z+MS0uHYZuobICGNmh+x+J9
9hroOxXBP1ek0xcACSnN9uhTV/k3QwbvxLbGypBa5uQ5jgzjb80gOF3yOnfgPuxvEwofB2agCsM2
tYof0GQZrKos6OZpq2czaGD6fbydlDLBTX2DmPPa0Ia+ccsTOu9eZYXC22vIwuAdWLCaNIpkcoj7
LpPV8y3Qb8wwKUOVKzBOA6bhNSF356bfMjaLmjMG5eUBowYZZ5IMuGw/m40YJbU1OQQHPoAol2xo
o/PdGm1siDXP5kIuicL60uy+ty/o8yrt+wFYvjNLKGr2Ritsxfgt/BR+/EOZRe1YLLHg0apNL7t5
ru9JBtM3C7WUkABrLx1Gqa2L96Dtzpn4gL3MGabK8Z+FGItE7L4fRb6UzcqgVy7wonAlJ6WvH28Q
H/CeU+GowkcocIHfhm8158LkqlqMR4MKQJSE+JmBJba88F7UHebmzAeX7U5HiiTJipv2HLJpvy6g
sSRykWy1XwbS+Z5mZLM1kbQkhtw6DhTk+HneRBvD6+r2VeNwSTmKktPC0dEYp70wTSJgSHTwbdeN
MlzEmbBL9fjmy+bYmNB2rt8zwk6V2+NB2tpeqNjdkTs+kQ7Zpvgl73ht5mXnzpdbsN5KtO3GfhSd
TxRreA8Tb26Js+KlCmOxA8rHRtYD2wWyliyqrW8T8tPBovCUn5r4bdUsfaYs2hPV9pBNxeBgRUTL
6QHvtQ6XGMLVfmjdFbYHvzRDNMG+yRKT+Tf9zUeCvfR1LL9xW/plJOmXt41RxQxjcKU+4flygiK3
bT/7t7yhtxKiypNeUFKDKbpU7X2iR1+nEgKLyUIHRbgezAkGEYOFATs7zFT7FK5Wwjf5DEswmgU4
y3CHTqhXtInTCLy+d7kIiCGd59dO+Dg4ksm1HyaO+l3kbEoDzQkfqc9FQGG46/tg9RW4GStHjrok
4QLIcYCnPL35D80yGHl/xcCLG1r7bFXAge18Y1nYYmsAHgY/zqyUoswc7DxvJ36A2Fnu4P9yJGwE
oMnbSc1FHqi1Hii6rOZcsr/x0s9CI3/zNaAT4KAvkO7lK/HiqiMbH0/OAxL+lRfMo/fhvr3VNLYw
IL6PM5QLH+axsXuMJqwdivvJqsFkH+1SNqQH0bD9jlLH4aGMAoIZ5nvdojD0mcqr5IZDWtNMiynK
actnxbbwOMPg5WgwlYioXPImruQua9nD0nTUvYpsmW/RUTNKUwGHVVI4EvBH5+F9xxdgMg/artN9
eNI3Mz0UvW9nlj/VwUtDLeEy8DxVO0b3WJ53wjhnpZTM+//LTdZBFO56SvJl8EzWuwg5Fe7PY1si
ixNJtPTtEIDtMqH1whKrpPiKfc77OFhbPaNZIkhhNe1Wih0/+V/QF6eR6KGQuHaHvuhStuuz8DPz
VhU/19REBjux8k0sRILi4f2tKzwypbVSk6zfUWnukM2mfxTT6vWDBHaFGVtEE+PEDA9XdpJl7esL
I9eaOOxy4P3IluvUOXAGp+2GMBrp/Hd50Aq6Wy/kSpW3/rSu/luWoCDVhiEEvEYeha4MVKBQDDIn
IhTtD3nSgGeds7dwHvMbe9SUGtt7EjhdsqoNgsUHJjCif6WKG1g6MiphkR5T36wXVbmH9u8jAou+
JHgP+6Jd5a1XCs40q9jj4b440UmTIY6xK3iKki4TI2hJdO64Xg6qtDD99agg+TXE02j7lFkpOYki
k75RdECORi5nKx4L5I68OWb/76c0ebPTqrNU9FNPb7StQf/pk9weMMVfaUp/e703xpST+7BPKhbz
PKDFqs658n7z5YoExMzPSi4YxwCod4PRqOyRF+xKwrTwxu9AfGwgj3lGvlO7v9u2A12PvjS50oEx
jL03AWhniqQ74pK4m9M/kkzgn/4DuP8wQ3Vic9g0qBYted7ABYpWxka+CbXVIz5mcJl8gAMfURKA
D9Vxchm4ekm13Zxg6t1wIdDxXB4FtO9usXFzuMYEQXoNoV4uqxx6Ua8yS4QR5G3VWGD7yiSjNK1M
9pNd4zPemRQV/sdLlSpQ7to5PZWhex9nz+pxGtcoawZwdOtBfZ8hGu4SL7Cwu6yet3aDLavHgcre
vxHIcMzwx5rf33fSpEvs1jjkdWwLVU/sISgPOY+c9U7IVhvzxujOgSNy/kQ76dE1vFM5NFU1k4c+
tMF/ijrAPVSq2XKmMCZdU5Bif1AjljuOGRwWu3rs5nLUmbSlUEIRqTPM+2x1iWCR4SvBvEgdltlD
ZfNDRdWHY8kcqkv/MpeCnxgTU8uUly4//wJJlMeiRb9GL4lzeSGkk4v0holWQq3JUlQtdGrr9PTx
j2mtAT9FmUkA9iRz6Jlk+kU9hA2UX4fDGlSHkJc8Tj4vbozpgp3y6q8+HjPZ+Abv8aI1XtRtx66g
OkTyD0v7LnD6sgjPx5VIvCMdgkTovChGxSTlowzWGPKiczom/BVIxat6rbBpn+JmCtEVzN7+vZp8
pmCXo3Ec3BduUpifG7l9HviDxV/dSP8qFXW8UY1s102CceLB7lE+hmCtyMVKzK+M+WkYzkjozTUQ
TvKqfxeYvtGL5nDwC2a+RvsLQ2z9Bjusy4qntFfh4PlUYs79XDHp3Vcyr2O06EwT29QkMiSZ+zxx
aUd5MLJehSVsZJA/LVdBs9LJRGC43khONJ8FG5YtmK0ImojVvMfph6jDEbwRZNwwOtnWPGAafTcc
gbUuDnhTM+w4KgtJ21cxsaAAxPebMZETlLPkmd89BY5fWQ5sZ/AvhFDtnHp16pid3cykwBp6ipGN
wCKszaA2s9T12bUNTQMUAcaUN0jyr59kRH20gHzDqqFY5t+waYmlfxVP0VB79LAntJ+FryIiwiyb
FqIMNm7HZrfylOkL6EltfJ2OVB5DqQJb7TY2p4lXMjSsvKZjK2qY7NEBZ9WnrFjiPka9hEEvfxly
QKjzdCUcujAgSpheiHYt+nejoDLTCw5AhE/CWvKDoleWifxUdojHX7t8zelVvl11eLb4Slo+LBbQ
lpULjfmUrLE/d5t2/dui7AzYUiEvzK7kK14Z2RjTGQusKe7mdWmqTAHtGF33KF9gGUoYF/pdlHCq
cLPzKlJybt5zvbdO6PmPF7UJomxwdVENN2IRAu3umtg7fXrMDWz7V6EU2myD/zDGLAO6uLxgsT9k
B+spSSvJava+P+V0fQyGmm4QdHT5xymwYjjXXA61DfdsuJSfiYBHxx2kB9pUyKjFcgUzZmLARIsb
ZoP+S/FrQ8Db4hSkepQfYeydcgXL/r0YFys8U4NW9sQlu2iT7KzjLLIeKmJnBnEqwfVzUheeW+/5
bfK1ravPUlGeu/iAk33iQXHFE+iEY8fvBVNlMe1n/XEFFxbneDaUvDr2ayzt/yKDRODXpFp7tYlc
VSPqj5zdnO2IDM9vUx+SRFr5KGLTdreOz5JImdQOnmNgJqz5G1Qt/6I9SzNCec58SU9CUe1jiq0Q
AJmWPR9FLsOitbUIS2aZ3PVEIuOg04DQy8E29p/Esc5UAwEPJ7W/eek+3oHeqBKmlN5pX/pCxm69
9sFNJw7UZ6DeEkKTgGRqZMaJxBksMT4XtX+GnbvHoueme/J8mrGaH/sP0oMcyw8fg1KpGItYo65+
tX8XrW3/fkrD61DifubFiEeW58fOdCTwOD3JrjwzcTppz+sdimFshmbA6WKwJhOeZ+cxQVEVresK
oP6lZeH6qAcL+Sf3ET4e/klA3edwIMusHKxQWcCJPm+LIw5VjAmQlNHW4UbXMC2BokWfOtd6b8go
2xfnjf8s+y54KuAwC8ATFKtvR0UuLvE6VfQjGFv3jCefx2zdfPLKy2eV78YFkOnr94Q4ferLeDQx
TRgajKAcFY7J09WtdZAfo9dV4hFyro1yPltU05cl6Iz49tf3ePvIA1g+oY+atVkASZOeARM8OAPD
+Xvk+2wWituySE0t19qVS5sAOQgD0hDqypE8gmajM+yh140m1l85wJD9nT2wZF4ArsEIokKe9P8L
iX/DqESnxCbGOq5NVoq2GhdSdBSBoVdm+ENVBT6jRkKZsxfDI/2Vb8Gb16bTOaIO27bT4FKeqNeU
3IOyjaL0WNzl//BBCNKCEl3YeRRBM/X/KTHoWUUzH3fgSGSsEGVdE15HgtIrFIiaHo5zbAVncHvZ
wGHnRi+o1TgWYacrpWyeaiz4dRu8KW+K/VTSE34bh7iakO0srE/GlwgW9unOXb/FSjiEb7T3y2IQ
lXuXfnIXSK4dgtuCUeGw77ir8VfVpRYVdDc/jyBvvlGr+OCAiIZEOd8RnaLtaKWMDgWutVriOpqB
CbJxtsfhv9gc+qnKOdy3vu46RDDOyi5wgAjBLmhHG20V9frP1Bi9X7QhwJIaMR65n2yEir/Vg9W7
BB1Smi8oksNsCGA4tXnSAsNsQae05NpHCwPedxVxjIrhO2/1tryTuM0Km7DmRqluRIjhYP0fRIXY
8Ij6JCEPbuAUxHAeyw21/8LQw5CHXFWIRcgxV5Cl57SLMDAGyzWri/AWH3OvRNi/i2gjm1XCB3/B
lDNB08z14q0MdEUOrRwpJMo1zLpz774IGKsp+0ySOt7O8yud/5OH0OpU/cEcILVuKPc6r2Xbe7Yl
s5iLnwYkBbVxNT8TJAmHyaJsvpuDIHWs1AqkgRQ5f+nvE4oZu2OSdtOh3WZO0xsHqLWDmqGuM/5E
q+MYjH/Hj/r2IXKj/Idlv1V9a6yIf9TOezRA+Nfbh6fq4R+8LkNNJcHWC3xz0nklUqKjh/VvrO2q
48XdqTgz7vBLADu5O2PKUgacMj8ozxIBQz1AOx8hJNUCWk2jkjdhHhuAkR1DzTLc7R1D44FPvlxq
k3BXkUkudmF7g4XXl3ahbpAHqTBAlp2tbHmZYMM8CT2ld6rE9ENi0PWt1Z1fPMm77kfGGgp1eF6s
fp/fzhBP+OSV5044kz3CEjf4gKBynzdT4UM+UhFs1r9+6LOFzeoGxItZMgnYWMNCD+CVjgcXo9a0
x4DxV4ZMDwgKPHycn1rwM90aTrDcrYX/vEosp8g/rgZ5Xr0wXPa7XZQcfsTOMqhfCmwkgccbmO/V
AQaeC2NBLrisYgcBcuEGSl+nLBL5o4CnGgHq/zqDwBulq+rEsaOPxqRdwbGypuXQsKoaWfDauIzu
HhBM8tf77SO15WHurawX7h4nK687kAsbbikEZrnA7fvk6hw+TeMs8n1etDROzr2rgZIfrWRE094G
/9XXBLJAOquYj6zb/zPt6RHd6Zn+cnvscAuf2M1UqjxnzyQL52cF+0TKTPA8uWYtn01/261JRXCS
OPxerZvsPlVCWWkmA1FFjJmzKkmFZpfWKoaHV+9qUfoF/LkrhU+dqfHeUIjJ1hHpCW+vAlYKH/Yw
mGUZ6LF2HDeSCPSmuz1LGSQ65nrcQniuHSXLGcVzoJkDVBb9HCrk1cH9fn5D13EUb0twaZEGB8uh
umTtskmkvUgMd1j9Ztl3DLdZEXfY3CMTOMAr8W9hXVYUkjNj0hPXjel8IqOh3cDUSzaEQvatc81Y
MLNBRrW1T/q6XEHw7H8An2LK7JMdScpZKC3Rh42swFoI3K+61Ge90RXHwuDr1lOdwfMj1dhoL03P
9LKSfxAQ2hpjbtiI4Hl5gRIIIJhBv+v9C9dEYYyywZVKg0OEeWlzyR1LCaY+6KirXFqMF6G9Szu0
IfRshIUc4hIxkhS8gWIsQbyFWWNv2/5tGMUSmlxSb05PWt5S90agK53fDDU68bmOidZC3C+YXIeD
4Sgcu2rl9cYk4BA8rjVaiwzZ+PnozSFs/Uy3J4JLPo7q/Lfd1tGrR0tO8WfCe1gm94bKPloZWT53
EDpx1X71qtaaovuU8lIB0ShK5noL5sgGtxYELCQBst1MmJjh8yG1CIxS4SqOAwmuPF+VRQS5Hhb9
sPf8z1K6UuE0DyUSRvNjv77c+4/v7bI0BSqkgviN7gVkmH75SwZaW6tde62xAsnHnVfV7KI4XCGC
WJjZkQL+rGYqs67CnvIl3bdZvsbu9LUVL7gkA4waCUa2xuSuU4MkUFQ9wk0cBZ9yGMGUM5plr26X
rARCzmzAKLvnp39N7k4ZjaCkcFIgD5IqlT/HTcK2stdOmbI+18avG2gUTQeR7Y/VBXFbT3XIuVOB
uvW0X8IIj2M2WAa1FP31TQ5vlDTamIiiGc7YQj0JICHp03R4O+nw+WltjdepqKTIvffGSTqFVk2T
HYdqp9qcFdAiTd5QMT5hzmqN5hCdHtiEl9ue69vpE1DUiBnfsgQNi7KBcuewnIKjLyXapKVr2GfJ
wgo9XMVQag5qsonZx3IFrfQZHsoRD2ADmSsZTxiSp35sheY3wovBtWgBSEklNIe50iFaHpuYQI7t
JaCGBKnHMGb/NHbrqeSmwHdKDeJyrO38fYQY9vV6zBFv3bnUvOga09a11xNrQoO6xk2d0WPwNHq7
cYICISl/Pd6U0KQiaIdbawUpmjBITpfzaw01msVTCGGzoo7pCUeHPiWVpoaNxJIwWqbbHWqxNchV
1qsYN5wQoLcSDv/n5wVESjdTm6ck4OaXxhQFB6NY1eeQMiyhJXhsr7jMo2GDmmSKRfmqWkNmx6SJ
xHKpFZBjzlvs2X2wOGnnr7IqMFG/1CeBLFqz9cZlMXwG8mTpFgCiyXyI0/AryoV9N2NIaKy8m54q
Xo/tkIEra3GuN9OYm7s+XEuLNJcRybAEnoLVy5RBGMZRqCG2fWRXjYo9NxyuEjL/SPdVpVtPKCG/
tcYcXmpkaJw2bAbzx9svhjoMSjnvNrtMXJFu1JwK5o64ZHOi9Ca2O4/qh65aL8VfsrWlNEafC5S3
fx+EtESh490CGYQ2fWj2nztvSYNLWLESLElWd0xfqO10OZ2CuX1b9jvhmQvUj0CAn3OddsIRiFKl
TgtR91BMu+x+c0aFUhH4KfYQzEzFfwK/8w8ctxe6gerfdPSyagSjv2qWZDAjNCTFpMY1TT21ZNpe
CaEK315Qq6mcBeYnzIo333fivzY5k2YqkaW3ERpB1+BNnDMG+w1jJce6XdmJr8cFLFG9LNvwhCzl
2YO76uoNIv71BdgQ/SU+ScuUMcr4B9LVadQS32kU1+6Cc1U5oS1zIRIvqtKmSHFE2wMPery0kDL5
HDpLt/V09KUrZftQyqa7zKvUhwvRriZnMe+WCRAIqECkmnp4XqCOTmbMYwBjPYgWN+8n7YgU8YdZ
cbIn8626WdIq5crb/PQHWX9pLKAV6zzgxKrVwiPuFufOjaJGOjsgMVVRNXx3mxQz3YTK+Uyuzg7u
2Gom4efFVX0yhBV7gDBz/0lguCqU4JBH0eWarqxvIIMaEQ8TI7UY9JFEIbFLCHYbxwUCkxF/Fa+k
j00jsnbMPIBU52QWeixRkao6SCKv+ivOiomUNsKd8mL9U1+U0MoXtthevxbbqPw4WqbvC+lXB82y
ZxBmTFCPLXZrp2qxpBA9UJEjKQI0Rp/0q/31y1XkkHLfx1YxoYkPnpuM0B8SJoh1UKbvDYaAdJqn
yYREPXT8Az/ZnYrS7qR9fFIxrANttfiQ70N5NDundOnaQe0hng4gj5e7dJ7b9Eop16XIkBKG+6E7
AGfe5SORO3poaPAPuhtnGBJupeZc4Aii1+peZxGULHMwEHE1/X2JJ3Jro4CA5wxlk64TgAm7Z+w3
Y5foh9n8n3SAeYhCp6cCjQm4blcgHfs0smTVtZl1DIY/L35PlCDfQxnriImEuGqA+OB3u3kf+kWU
sL0IK0Q3KxkcTiZYYr8dnLOkRonbb32ntCMdyEym8NT0anqRFqGFl/5odKEUKwUZMVbYGKPgwQIa
Kc+8Z3JBUnXaeBbLTeN4ys922DHM4YzALEpT6TBDP5TVTuqoAwOGKflGfo57w0c+yfNQ0xPsmrc8
GjqrWJ1GKS1Wa+Z/Bw9J79lSctmpOsERpwPSxZAIfL1QbuFaRO+NLXSlFT5oG92ANhAu8aKhFPOE
vy8YsNWkBisXA639L24N94xCBVw05ygPu9z0mF02hsEx3UCynr4vO8M/SQc9YjpQ2PsIZzyeKg73
DG/DP1DqJVm2chCHKUsiANDnFS2Z8q0VqsrtGRk+Eg7JVgoDtkaK2Y+hulFehaRynDGei/skeqDu
sK0Rbn8AvrispTozvFolbCfIv0CPOQFE0tdZCXklW57cmddIlTAk/zo15nnFwL3vBU1M030VAGYX
124kZ4aUpQ5BeMe1EkMbnQL7h81zPx4ADqGrdBW7x7+o2+KCgvHftbENolfP1UB2zRtSV7x3SbnE
g09/UBOzKwcP0mfQVxYRtZ4RFe4Q5+6BI5WCvBfGk7Ro+FuHnsZP2OLyyOFxGQSMI/q1rfLVlcLG
AHcdNrLD255u/pJm3B58m93k7HGRI/v6RXYd32z1yUrty5aPGcN4FUhENHG9CYx1Uegym7uiExnA
RfYCOEB+9hp0BRZThMkfMQpjEbKp7D73ZDg85pxDtBemXpPr06l5n0tliOrx5u9vCtzlazAEtM9B
Adak+nmSZcp2WAJqjHVUP29CJbxXuaH+BwwEdZ8+1oe2+X0bMP51JaCDUmMIWG+nw5UqHuX3YQL/
bQz66Rb7UqTP6B6XqR5Lmp1wBKNRF7HQQX7koPnhEQ0L/x7jQLREDznBXQiBlIfEirPyf4bkyqpL
5/K4JtRavlPiHCiud9gyAG2NpZ9+/lPb6nppnvEpf/QyPczkZsSasy2QpKT+naQDP1asjAxkESrl
+vWoo7/QucXHblGcR2E1At1dux/AGNdFmixHE/P/tmrl7p1R8YSfsq4Kb/+QvcKQdPNwr2ucOBxu
qJ/WmV1QiNNqEoSstKQIdTj9xn1q5ZVqzwjwUWcmyEpmDJ6x2+0efCWN1n8XdRs6oxH6B0jWave6
dY8gRNnu3Kaq8Sn3sCjAnpcOvhPQXze1BaOmXfBFSE1pHNBQz0NwcrIGjg4NzUqpnFVUuCh5cGEe
lwydpu9h7y8JzWvR9/Fx5uId67jYAc1ayTPQn+nH2K3ZvyCWPKHSmLpmQJg3uwzuTcRePEQzYb0D
9fbs0HfnV84kLtWNEAynTowdhWPt2/gFYE1sUSGEUGvXfP8YO+vMhsYiNUcsklXtxyHthVFydZQP
jQsnSd9+h6FAN5k4q/5DdMFyuX2qWd9ZFBxvpfUwxOIVdnlZPlQs7TSFjYFY3Y6fNfPH+MbFRmOW
cKb1vAj6FyDj7MV4a1HLjWLyvqmrhWCykw3LcsnpIetAdSSBju3X5DXQrXZ+jABNFpEDEc5ssodJ
NzXDiiGZVYrLceB8y0jfiXUKKM8zBu4eu5ABxNYgAk0x4aQf7DU6KX3uEAS7vyFCzZSXHPEBsBuH
5XNwzo89c7uHtaM/3CmpQMhiKhNNG6jy2xDfdGcO6eWcHU1LPEka/1Nh9FF2cNUr4oRPRABBH4K0
Lh77ROqznaI82IpdVMuWivWHx4uSd08zmaRPB58xSr60AW1ecxmNgl6QuSrl5LBOtV9eKF9VzQ1/
hj029rvNR8skq6kZOcR+S4m7QYQhdqb/dNOlVwTYi8anfHxOC5R3y6AOy6pr6SMYeWigWonDB34f
4WRsVulyj+beG4cvhaUGbIKW+H4ViZ9eEfPiMoPN9BlnmyWcnh4tzMfa2LFhsLze0a1YkyRK0Hk1
qFPjIGpLtbXMUJD97meTGDJlVXOnI/AvcQ4uVICevQy6PXJNwgOxzx2El1nqRwALsCKaMv+6tChb
UT9qKSqiMs/7glcxTAEy5UD14b6Xaon+0NY9OwlWN/FX3s3GCyCx3swHRb/BAa9w9wBXvxVhDRX6
IHmQHKbJNuDrigSJFZ2n/gF98onfwlufrsy0sUzYBbkhAnFjziKNEq43zJYut/iovBJWY+9Beeet
B+JeNOwa6zEIHEfbJLajmcfXYVGoCJSny+fySO+d1dW4k+BMgsb9EmMnhW9GKuj8R9myzlrL6z1P
ot0Q3/1jTF87vsITBaiUR+4NwOA5QcSxv8Ya21+qTyH6IDhjz3nZaN+delBDLLCY1Rdvm/sdKtvO
tJaQ5KviIuCEuC1fLlI34Yq3PVVthF8q39vQ4jNWA+pjUIPprZP7U+F+99/U6PVKFwAPBn6PiHWA
eFYgXK7lTo0Vedl99CUBO2I24Oc0lM9x2DKVK8xiREWzyKP6f7ArhVhnqYQNDw9aIRIRZUcnF+fq
df7eRc5gXtRF5Fh7WTngr//d/sae3C7mp+kFHjFMZljBXheb5cP8mYIp7sigiikn5uV8JrDlzWHv
bFYH69kp8TuBnoYRtUZ9NWaoJFvENQF4euU/v+H44mVeZjGoV+fl6XX1SG8WXfl8eSxRvUhDg2ub
LlDF8PGasHz3PT3e0DvhVGyJcRRH4SsLnaTbnKBMFgJE5s2dn1SVsoQIiTIgpzMOlY7EYRR4zO+Z
Wbp4G8bnu0TK5wWcBcI2hh3KI90zgdxbANqEUGVKdKC5dvGAFsXaQ0gCn99USYwLqAC6k4aI6y3E
ccQSmFAPfmXsURfWCLmndCvXC0iG/RaXaL4ORo5f1EZBCeCL1BA+AB99HeSeyAtj80apzKE6SEvl
g6qaLpdACDN3kF0iXAx/EUn+kQ/qPDTlRB/rZ8YViKr1jJC/LUeeW/ohAACntcJHxKDrjC4WZxUC
DRQfHMQhhHvsP2S4gCuOd7W+v5GTJjrgXSofaOcdGi45JctJ+5tFh/3MCzovVtL9KOfE9ufrV0p1
Nfbjz8cJ1AvtCbiD5taJaAAzEXpV2GEZpSq90gGqw0UwD+3whHF8NKwq6l9AsU/OCkeNDZDQAdMX
VF+25+tALFTIa5Z34pHVr4Q5gt/Mv9D8PhdlBX3hXnZAoCOKgEhJ7tXPNC06Jo1o/QdWDuUAjW6K
+1/8Yjy4ZE1NAkVAY0cIIu77MdlekKo9DgXCptF5WR5fcGQvIAUQ2toQntzTUvFuNvMeIPed89X3
NeGpA7c/fM6Mm343ZrMGDdwKkDeaXdi5REolvwceV9nvZKehMIa8hmD8wsPdEgJvUxGDHHP3JlEq
gk8CBxe/m5sbtFgvcv+io2prrVIcaD1Pvp2D/6TVw07QZfxotcU0a/ppzsuUVa1AkbY/O15f385u
/NZlS31RjTLrHbscrVTnblqQr9iTtOem5030VZ05PBvAkTvTlCEUWZaUcyErrakQCZtkGm91Y+V4
nKgd1KUmZ+TppHTd/beFit/DrAD4cEu+wWIKD8a0iZoyB1ao8/yficRkD0wUj85B8kRlBMkh2h36
DCp2LdyZnl2phiafSaPgFxchDd8hCHVSjA7jxg46IeV9iz4i93wBMrdXJwXRjCksTiedV1VFQ+mq
IcfFkDcvtn38VMFd67/+9jUvtCxSXu+6s6SLrOd+QUQcdUDihtYH1WaktD5cEJbxSx6Gtpe93GUz
3Z4X7x95GLVi0i8TVhXQazCGEliFxMSAnMlAmvgpfj42E79xB6qKrqfzM1r9rVmJWMrIDASuNzwv
3VYqzno2ffM1py7emOHuQcDQlalM8Z+W9gaIhXCjgMBtTSb4t98f5ZnzpNpOA2Sy1k0Nlz/pvOtu
Ypj8n4BVLbKaQ8g+JMzzCv/+az9iV5AZAhq6idzpcq3tkLQvudTnfNLpri5OCz29FowfOxa/8ZxZ
Ur8q9HhFaCG4L/63MFyaZDFo4IbiXhVlfs1iLA1g8+DrorAXRkRrkTWsWbkANMuvpfxNqNTvTN59
PSL3yQVZszjYoIFe83sfQQ18e7ttuNsRDhLSfLywYY7pFTDVQmjUYTs7NlBlszas2GJoBemybTF/
HArR1nQ6beV+Lh5LppEMrdaeO0wLCm0LslVDghqwx3KKSrDsEdFUjxCxneI3afuxJFo6hAHPB292
p04/Nk9wBW6CX0HsPHgPEvz5Y6z5DRYIObT3JwUkjmc82k+JOdxGl0VjQcFQO+brbTDASXlkJU7K
Klz5/BZltJVVUMO6cazlHW+917ntAEKG5P3rRuc/mISAQgBBowX7CMQpzSeSSrOGg7ztGQxe6Peh
vZVaqUwXmZlcFGNKx0yAp7c4xnvuVcb9/oswDpyN17/ypmjIz9KkMwarl5PgDbfIR1l8Rc3qJ3Lq
s5QKiblfmlPXo8ZqCYzYCFvCHrNqU1kD4AkIy+MzduhOTfZIXpaOPMFjgQKV/Wm4COYccwwo4aXN
IsL9aNm6foXDSlM2ACh/JPf9x8F/158xb8m2An+11UsiJhONuLMBguK7QGg69KM/f7MASl+5Lmi9
O82QWZzDEpmGoIXYjlKZpGA7vjT94RSfENxPKPyrdwcbvaBe45fp57qnGahCfqUm55FpesYc8kt0
B6ZMjAZYBdOIZ+niC9JVBX7rga6n05lt6w1AcmWxRL0h2Eau2cYsYKS4lnzjQFgVO+Fa+wXa8CGG
eRdmmKmonJMwWjyMdpOykuB/xm4qdB0P6d9QiWC+9u/BpfpvY7oDW+aY9S+WD6z7cWCU2NJI6hep
MaeC0vPiYynyFcBVx09xxed5SpZ7MnQsmPtrF7W8mfTlGrCnECYt6iVFordPLP1XXhPm5KkyJvqI
l9pzXENBVJnHTAie+T7BDu1hsxmvi3Z9Z1nB8n+gObB5jfbRw/TajpbCbDWrtHa88JQu7CuS2EuW
MHl6rYWcF6U5K2tm9t4do/PD9LYNaE3XVWq2KpdjDk13RQk85ydOrn9rJAT+0uTpgloTyfbGWr78
jJevlC4R4//rEYTLTCDHpPZpXUUGnX+O/9p9Dmy9lJwBYWu/Mnx896/zWyTvUY47CmJnQwJu8PJ0
zoMXWxqBgBZ9b/OYFWcMn4skM4D94KKHPX8BArhaUqqjYrs/HQl1wwgreTK4sYyV27HHn5NxSJtt
B3UfZUZ+wQ9tcSXLiTYMVgx9/mEnFF9CgjENjRxopj5UwCY43Ykee5KRLCP209wlhnC7DhXXcAne
M2HZqepQQDQxZX7bWK2tpaSoufm3eAk1DpsSXkGqaVqiR0WDfyssj+/5NaxE+QPVTzOlYisdsZvU
zb7VkfURati6ww+sOSJtW9H5AkrXyRKkw8rbvV2wbrPMEUWF7j103oECGHeSTlNQMHSBBCbLmFgT
A3q+nD+xMCXkPc3M/zpdJf1eaE/mBl5qGSsjnFntVgIAw3jD9CgVtswYn6YZMgcLwWx05Ez07JbV
wNEdx+cBN8kMdfclpF+RGScNCBbmeGMloPt2dx8w9XRDj27lpMMeMJu+9VxsZZHe19Ge4bMJqtnS
EakbgqLJ5ON4o8UoZ4K5elSGTsGBqZBl5qKbGeqCkwfs1dgPG5wBzcgCVCRjGgtnjKeyTIDdjTlU
l5SoUCjIwQH7suhUV0s/p37P1dF3FrILfpz8kNhzKncewf9O2vWJuJVLP/OjCo6zefTMAogQwAWd
fCkFt1NPicgcedGc9CBrTqqUd83WFehsu+iHJY2XKcrrAStoZ8kyjDQLf6n0HbWAGiV16pPVlnk9
OzEa01/U/9zyAqEBAGDruaNfft2B1VF3a+1809gcFWM7SIv6rxfC3Uxpda5AA3/6AL3uIW0kC5xW
kxs2KxYLchksm6Kpke2wsbLmGuUWF4vDMze9FcnuPU5bmtmcWhJnlhoZvrX7UxCr2yNpTOHPDUGH
0yl90VAPTrqEdJExJ42wh6Wue1Cmo7Vt7M1rrI2/0bxoXuFOOTQsYZy2yEVN8MumiQ0Pmz/YyUR8
QIM44K3o9O0ho1smqJbn4ab8LwMT9B9WyAXLtjxGI1Mh8HiiBgelELi+SorMJgLvSjkOfY99tfOD
gcdGLdmpm7s+1V1xYQZ4zAH1lhV+Iy/1fqOZoyoYklExf9Sb2IbAcSCN5BThjCZz5mEgewoDS095
yxpBLKqvayClTx91RSGLDK22QVbsF0ahwi9pd1ktsxO4zksQhURfW2Er4r9oMsgx6ni9ISBeMp+/
vQhjySLR6DfuEqSDALV8+CkRgVZaBbMtkCpk4pllEqA4VNWESpXgopV0LOjbCViGbZB/Pev0DgYe
mCWRptcW4YvrBSo2o+xJTZuAciwv2WJnXtXbFFPlYCU66yFq4QwI7YMEUWYQmMvgW7m2KKh4rpyV
fInk4Po4RjeAs9pZepZwV7MQKM6XcmwO1VRn46fEKWOJxLzHSbeX3mBCrgIrZ0pppfLmtbHBS4Mm
bVD0WJiRHrgF3izYrNtrdtyTsg4PWW3TOCOjUYAgCBhOaCAZKNRQoUlWVbmqfuAyqtuwdnOoBQxh
w5zRLmnPn0zrPAmuhXv8zpnmFDqmjvK9js6NcyrNXKYkErYuL8l+G0NWkAyKKNJF2ZDZ0UwSRx/K
+ytWiCCq/hxsW1ljtl2Nuifu33niqL6YheOh7q+YXac5Wdw5BNBanlkvOMeHzVZj6fAM6vnseyOE
ZM//IFgNeX76n9dPyt5M/UxMORdCeqcYoCHS9+V8Z3ZgTeKzlJRG3dTWJ+iAUaJIrQl5sAMpDNnZ
IiF2+wIvbJPNVEkJQS9pppsDlTT7ZCRGqTF4smRvZ3ybS+brKWxe+HvGt1P1xz33Csjj+t+fx0pz
LX8IwLiU7k6Dbun1uSPl+C2bggRckijZxWdxndAeYOH8IGfCCEda5PEC7iIBmnrs94ov+/JuGu4c
LlBgIb4P7BOShyoF8x18B2Wo/1i9NbqC34lqYWXsFGGx/7sIy9WWO9O+y0aEUi/mCWtTyFEtMvlZ
+tIAfSMfh52uVO5fZIpi/k0ubjLtSDur3bYJIJBDFphn+gaLdzGWOlSSbLh1zgeg2nQt3UEfqJ7g
31it2BPA0rKkyGDiim6PHwGyJ+atMBihPWNhNQNkOYaduZf/RXcmcxZcavjgqCMZRBdiEbmpWZPa
UBpWR5uPY+OJSR/KLBuN94LtobJ5UAr6caxwFL49lscWXzBhZi88q8QAyO6Hhn1BcA1O5YGnD5qg
Kx8nfb9IGZbEVVmcsezJGR1kRfjr87BobW76LuNT8cpl1xBX3PxRynkCEt2AJ8K06sIBvuWAwqTX
1kry3Vd0iAd3o+17iLIssKLa0MWI9Z79pXFzlj5CEqfDe26qpWTIDuR326h0bzIVyrbPcMtVxVvY
Uq+BDoNa6q7UPkNP4MlS9UNQ5apkoF3m3+C0Npt2+T59Env/mC24EXiHu7/svf6WN1eB8G6FowKC
DRXkvXREb+M5DVKzs7fhfNuCdsgYX5mHRvUJ5gKBBom7XKX3ZE/Bx5DxnDPZmtPDt2pHR7q1LvHn
2ZZ7brjkjRcui7ogYPR2KPLzGV7Bh+gTe1ZEwXEFNVy5iajl4UqDmi1qpYqhaCO1CuuRokH3m11x
Dy50b0bLY4rEFT4/IV8llRSCmmtBDIR09zLts21YA108Jx0T/r2jUUtMQSPssERoqP6JzxlilV0p
7bJ2NnQHuNgdzCNu5S4sl4SquUL5KDvjsuVQsDX0hfmFUMUWbKBRlIYadR57/qheNjlAq6nDPBac
zidkVmtQtxupxRhC5y3w7ha7yttJHfRJx193ztmzmMn8uCUYmqpwVgzfMAKFUqADvzCXmkAONwk6
n+u4lpqhQ5udFBOtV5fulFD6TrCi6gitfdT+Ebrz0sxHFSavVk5KEOMis7A3vOqnV5c6khZecty9
gnpFA3KSgFDnzwnOn50qLB+N/jCczNeA+raXYa3Iftor2V8CClr8sCQC7pQrzUHNfxTKMAU4ysZl
e33NCzig57fkI9HA0nRtHBMiUzk/QFMyE/AizDTiMt/yNfFktMpv+r99CzydWT31t6yaIs5Phu5E
kqRA4AmFVyOMcNrrOC+JtITN/iWnEB2rWuvkYJPcKVxVo+q3wtc74pzaCcx07kTM12wWMePj8qtp
t6+yj65IA2R1lIcDEVaaMP6EzJblqPDM3uV/gYllzV+m4FoQ6acj3Op2goYXwAvYXbvkmy8fRpRP
HKP9yfLo+CazmbAUlVQCqOrPJ966+hlTypq2y4c6o3Lf84ifjBfvCODGRszLAbn5gI/voAffdjiJ
DgaxSzTULnjIbcGWPPxtbfr3ML2lKFxHS4fFH8WqidlH9C7NIqWYH+LoN0o462+IkvMJA0HaR7G/
wNYexUGPX8qhJQTaqHmVvh7Em0ufXKbcVSrT+Nc7kvhQDuI5U3lbrHLOQAfeDtxR5u/CPOcfDJQM
zph4v8UMWMqr8/QKBV87LRGXDhf+tXwdHsi2GZCUBbXEfuFqopaoZLT1aAEpcX8GMRzy3UzXTpJp
/d3GvI5ZnT6t/juKCfKGp+PjtV7cGhHVj6RfuAr8OgsSL9/vtmmn+PjOFjpucZrP7ChcTD2s4jMZ
dgzlK76szuGjhMC+nXXhO2jEptuA235/2VREooFEz9/niNGTaDpLt1TfFiHsSxzvKrgLVnKzzU/5
4ZJg+1HZUezCQWyEfBvqA6h6lvhwxavtUtmvjvxDtm0B2aPH5uk4+7h5s9i2NEVk4z85JSamhdCW
khVohMBsazG/7PiwhPyiIpehjAkVDVM+YsnYI7akcN9BBTROKgFmXMtQ5/C5ya/Idqk3K9keQK5n
UZcreWsoII7WN0LbtgybrDTUv99ce/2gL0ZSWplUFtyMjIqfo3LsDCbMvOn3g85M7AcbM0Y3Kk7l
issXWyb22w5+6DnCtqbz2/zgCMVi9x8CAOu5jGmXuCvfAeX7rH9jBgtezD04j0FjUYBpPWBeVAkl
JI6XDLuk4H0xSZImcgObmkj1OgVXN44Yr2QyqmAzSuhKKeJ8JQ80g9n8oNURW9POjQMQNmQXlCsz
Fkuih6VBRr/tqvBtC3+9okJWehLZ3O3vNfxEKJo2gvRTNKgc6HfXupT2Froby1gWyi91SNA6yUdK
b9lHhFPBg03BMbBoALrggtG2soNYR7ibS4r9IBkqHp0GhEHnO7lNZfFkYduk57svAgdtp5s7zBZl
HNKjYmKa2/fRHObYrcLqCBjvJenVy+8cMnFNqfSUlXxcLZJhIljlO8N9nEdw9RM2M+edn2+pjWOI
3eJmSnMbAG8KtQa/9vW90GfQJnCDhBvznfxpf4xqA2PWK7Q5XBHs1vrRCRqsImogNoprsIGWBG3y
V/Z8fRMQBzokRVIY6WHrFUGjQnKTwvyjSRcETcwYVjPATuRipcOAazf2J8H0Akq6UaL8WyUecbQQ
cA79Q3nY/Sl1iBd4l1AwR3XcfLJdBp0EDG6s9ezubaucFLQxtoZA5aWQ5zWBH3B3lXdQHfbzh8nY
5cz9Rnpb0S/RyD8v7OctRisZ+5BTuGU2pW2d3Es0UK4d0eMpazYrzEjapGMA7GOh9KF+COuD7xbV
P4lH9nZezxY/OgK3p0fnjkv/7n1ABcH0qjp0nedeYJl3FZEZwTHOadoCL+1bAhdMtDTm5umpkkPZ
72/8LeblWqEHa4PWhmH63mfGIoHeZgNJK9iYF4JkkK2r98G938rWDqgrkDRe/9awyIwBG+m8mc8P
AyRchFmHxtSLE3H/XblF3P8Is0nIPIN18VJk720Ip3icOld6Zoz7LLhJiWQMopCwTikjop7fB1qz
AlbK7hbgKNr86hVs3DsSYpi98TntdHyvDiiNR0GQB70xig4GDWTyKES9F4np5VGORLpNs5JiBBj5
vUhR49/T+ilV/K3Hv9JKGislHrWC/SxKwLsQeXxdLGnPY/tj7PJufZxxYRTft5QOKSQDUd874jMA
caf4k818R9TIHsM7HnM/GIYBOkzamcju4jkeBvYktZFqS57GFComXfoZMwoXuFKPyrEU1h/FmxzT
eZiTq5KvyAVf6KOxupOFtboC8vewVu1+SdgCJhtIsHEup75yuGhRe0TassGx/Mn/8rgCZNZuqODb
8+SEa2OCjgz2CkkmzqnxEhJ51mbLWz8sLmNG9T6PSUO5Fp3K7gkMUYdq83km7eB6yAe/wq1WeCu8
20ttlIq0stESH12L1IL7KhObanBTxZ+U8pwidkMRKs1KrOeNzmWVdV0ZckDODNxEyY10zJgXRMwf
TkcdftghMVA7VyJCLH637HWCdKtgHPWdJ27UBi/NaYqSRVrqBNHME5fIglbi9x7jkei8tR8Pk0q/
3h06Ky2fXs7J+2JfObWEKELcCLJz8WGrBuQd6WUeoGKE053F6hQVWGA79kyodrjGrJVkxvb/hNZt
2JUoRqSFCHPMzJYwO5Eg4oZWxp/BwIEcrgEUBwaFwpHQ04T0msnCudqPfn2Q2suz5lKLdZ5DCcMz
OUbxhfsCQ433tis008ZaBwoP9uRGw6xukGFxKTzcZxa+cCKhiSX6XFrQpSsJvmAXhoFcumdlsGSi
yF188lCbI/NH0PbaPJJKoH6Y98sb6PDvlxN24vmn1PFnJSEpda/6JOvVAB3KoAwpHmMI7O6rerPa
bEGU7R4GeI6P09gymvJsBUI5UjmFeGPgd27OnxX0GI8l3WSaKLkc/83aO2Q0NVReftKnNyrkrIXz
tacm14olqp7w31QVt9gtPIwitMOz1jVJJgp8bcSUIlHamhuieu9fYgwWx3RjGnlmDY0QH0kguFX7
KHvB9ZcvZHRnLScbwPjNGdW7ziZDK73wChM9QC8gU29g6Gdhx6DECBEJSaeOcvsW6+k0Lm9vBZBJ
BcWWCjHFl8VvTSi46P+7y28ChfOQHpGNJMDzPNpz9x0zds9xVW0Z21Mc4stedjk7ghKyfUb1D7Wz
5QaiqTsca464O1UNLoUeW3V+kamiaCUCsGdgyQuvTwfOuWCvPcBu5leBbBRsyXIf2JVnSTJmqY1y
2eZG2KmiF/G6LQ11Cvf4AxwuGgUiftaliqkuE/jca0Tg6ZxQvRBczug6cVMQT94eEnrBZtHtXw9c
ln7ne/AR0ngD5XbM38TAvzOqY8aPU4/9VxRvSdCGoLac0/rfzoVi+1czmVrmLjU6jTxNvmv0WG1K
fh+klsvUdqEwB16gZl2sqzGaZRUzBC+PS7hAb4+WSug96Wt5rgIpbg6XskVka56COyrBs64y/2Nf
92YoVab5yCVmrJDgIg9zl/Bvb+uQI8kY0Y7ReAMWjrgikBYD8IWZCr/+BnAxRwukSUQyy+oX3oDl
6w/3gTSoXbmKuUVxAk3kEJAKAhoThp0MUkbhxtkAEYiJlNuhglVoDyO8OPPp5+ZRlKMj2IVLzZyV
EZppmeg8d8ltfzhzU0anbe6APEJOdV1VFKdB5RiKapxqu3w4WiMqUGyD0JC3d3pJ4r/US646O6uK
znqqvNIyLdTDy8xpD5K1foorIBj6OJBZFgHZGjtts5J642zFJyiNoWO8KV7kFRYplJgTUGJI9Jhi
LHMgBaDgtcVGWV85KjtoE7yMGUcexdAbJ3LsCczzsVYD1LpJtHTdnh/i9nVof5r4fIMLL4pehJSV
e05ZXaKulBODjWjy5E1sxSIRycoyTya+Q4CoClB4X5FVdseLRhIsbE5nDJQPuY8889pECzda57x3
oorQH5A93ARgIxypColvtsF9oTUEJC8X0PmtMgQeUDgSOPDK1ocSrNRkMpRhYuE4nZcjCPflWsTI
66vmOUMdYqkbrCt1nkFKoY3L2npoTUNGzBoDEw0PsL/2QbrIW/VQcGMYSretMYzN8eOHknXaVyV9
xgkqdbiJ/tyctfhertYNyx2/vU49RGQAlg/ydB9b1ZTTXNnzKV5vNNJ6MdDQ6TwUi1U89zonJh9+
/p64iR7STZT5AclEuRT8ZPgdQVnCMEolfCBbi+RO3Y2ZJ1lXWTZE7VE9RLNGbG+RBCX8z08SVXwu
/ynftPmxN5ICcEvKiuA7RdxoPdCPgPeJW7Gj2Ig6G1rHf8m8hsYNykIZbrivFHPgCWoARlaNuWh9
svjvBDC/29FSQrOy0vuCEwP5jm7K6EFeu7Nm4Up82H+hxgj+gxzWs9Z5oQxHu1w+DL3qYcdR1dpZ
JMR43JmKjwp64M0Vh+YmH6jdnjEYzaxXc3mCZeifkUv1nBylksPmWcxcY3MJZgSbw1tm5ZOBIe7L
JI0SzU9fyO3fELXKjYfQdjy8im6aJ3nsorBMxbe8BUAa5GZOioPcoifhr6QWoiSsLPh6XH/ouHPc
U+uBY8jiFa1r24mXLVlxl1+C4KEGTpYqi1YzSA6ArD53pJtSuNhz0KLsX7gjrKquk2WLh5/zNWaY
744EUmet6ZMY/q9T0gmJ1Wz6pND6BSGPDN6W/OHH088uX7phmzlyM2Uwev5mT/FNJsbBjWR0yan0
5JWpDqV1xJZN2BLqA2yn/i+GJk6dMjPD/mCGFEtVsflpVBHXP+8m+emDSpJK5Ur6oyBmW9stcZR2
OXchxX86F/lyte1L1w3yNxoFmcQhOTD3dzr4rrc3FRnWxRQ8lGNov8KgBEyqZaFrBKhRu8+gOFhv
Fh1xnQ+eHOyKM6bENhbE1TqeDKMkJLMOt4lo+6BcV64NymuCMGEiMTGXaYa63W66tFeYzHSpFw90
gA1HJxotmCpEoW8mFJ1ujwkc2eQijx7rLlEDnEwhA/muM8R05YQ8IyDWHJI5JqR03J7hT3FFbxIS
mNd6DsxlHDSJk3BkWIo7sXqx/ISTQxJ5iYMDDzMxpS3KsG295i6DUTbj+MiDrmnRBGqMKkTCvcFr
+reLsBx5CqGDjmRt4DCrDwFO5Eshwczdd+trNKYln9YJ50TgJ7P7lpp8oTZzOV3GvY6GMEkladbA
tu7KaIvjqoreMTbNnWPbFtN2VLdQEEg/4/DKmUiYyzM7SLBe5mFTSeZz7GAgNqkfKDZCL+FXVL4C
yatoSsSoLWOLvfKu33T72FPJksKJPktJHfP2oU2MwpYTXoqKjECTqdCZ8+1mmGr4bKRXgF7/oOgy
UAytS3HP3Hu372grJvL9Tld4WNey/k33AQTRKNzHtclAQRga3TknZcJUEt0KWVHquCCG5nrZcZB2
2HsAK0kY09fqnwGdYlP39t8+GNlhP4UVYUOyYUkmAAD2cUp4+74xJr/eC7POUmTkbutqCw4b/jZd
quk0dYU0DcZ6m+OIqcQzxVu1AEXtGCd6sqFcYN7sZRg3tLvtE09PbjfkXIuZZh23leRS27HXm7RD
OI5oUC1xnKkJhnbPNkvziVLk3IjYNvAAwy0a/VmNMiarTtEL2QlQvl6fD1f+0HFga8Tj+87g1sOL
tL2a1WEwfbXp3btV0NvMclooWrw5xwk3pG6L6GDXXfJOye+It9N8qt/DUJ466B9hq3e7OPJq5DIJ
O+mQavQROEuA2VeA7W/hWVmD3YZtZO8KI9y9WJfNXE9Uu+aHhtebWiTwg5PIK8vLnE/A7+peXjJ+
WF84/9R8hsUtRieK3uqIVO+IVIrHbdU/qz+2uPEyh28fH0VI4Uhc/oMoA1+JcsBM4dUTn3gheoEr
spHaBeFs9WDJO/lzR/QMTrutP205VuihXkb1aOXy4MxsABDwg1kzKUM/oeeEIdD8g18t5RHtfJT5
XTS0isJxyjqENM5yLCRQsMxYidufFgaNPIka0bQRlpy0yFgf7rvoPSr7aQsMdZABsmbCEQTiCUSV
Ob2/qQTI2Bchu+9Ezg4ZNqGpFcVLqPMNCKwT6uLQPKqUEujTfd/9LqQekI8pq6KWoN1z+EDIWwYq
cFfAfKgRDBAiga5/aZAo5XJoUdK5tRUDXpDJ/c8LR0wrwNNyc81o8oRWcGsY9ID7D/rqh0LuWK7X
wOdTQhSkMuM8iQj4f8mlFNzN9dKtF7XbktOXV6YfUg+aFeFQCHdZv8Uzt2wLrtbuJQFDwW72dk8D
H3cgfMpkJT1h9SUH2VJCHwVCDB8N8VA1hU2w1ze85adLxvKCsq2wzc8k2tmNxfLEXAnKsVuDGT62
qzMR4pcu+STaAT8+7AeAK5HluctDlMSMFu+mGuBWVHcd2ozg3VIMy/MymTl7DEfrf/5nZ6FZabRB
2J3Pi9CyMMHD+NhwF9H/IA0KdCtk7aO2ZcUJigBoZ+obtL9ec4sNU9eJZjem3+/Sce/F/FtTC1EQ
PtC1jW+CmA5XtxIXqbPXNjAMb5bIautDdphLvxXZ0Bx3Yg5vLvlT/Q0XsIzHJgUnF4VWXfO0UZSf
+vUiYhrgN7m9UIvuvqOS3oOE9SDn76n8ACGoHVrlw3YHzqPfIrXAzNQOyJNKh763cRySyCb2oQ/5
1pjKU8WRVwLbqPO2XvPgAMJZCM5bI1d42PtPAJxasI6qSRuBmVniWHxdZ5cyRVw+tjZiv1/lV+gn
N3EZH1HxjQ0ISOxRIXoY6hOq0UWI+PD0XANtUd7h7VirO49cI6QdJBEwNpovyQkuw6xwkvACqcsE
iyZqDYEk4CPvZXFtFvCzMSWDsWPM6qELL4InPuzlqjVZFX1lEEy2m3THxdQ0qTs9hAMWR/tQ3AjI
tWa0cEaYCdlrY6c1wBtSnyH0QZOPEXepKE6w2BlM4W3wIfKpu3xc4aAWLJCM/Q+cqIAoN9kzKn/A
MNDJIf+6qehbXVs3jzYfd3eqx26IKToy2gYrqlmj15C1UwUyoXagJhkuq4ZUKWagKvqRnXw9hGX4
lKNzbPrdSSLFQH4hll9mry6AmoR+F2fyP/QbqHCeqSUA6ZGtPDVu9ueFJCk7zYIP5Rn0oW6iCE6n
2i4OKjSFqnCGknCmFRBqjs/M71Y9cmMJnJVrs6cX0Yhs2PA8dCnLQPxZKVeaT5wAEF6a4lBLaLsQ
6AyiDqUxjhKua1I/dQw2y2Ou6v4r2f5l8QjR3dYGzfuRDYEbCL7fYccMGN/I5ciz3hojyPbeOBrj
vbQE8gXsd92LKXWoIdZrPYaopesewjhL4iBXRGJ7ocV5eewzkMYBoqrfNT70z5g/B8gME6VwHghv
ZRcSXsp6365+1vQgJKaABcYq9096CW5q4zzWZwXa2dadfd6U01ft+y34MsM1CaAW6d29Adw1Vbcd
vjR22Rie0s2XFMZRUEPx6A1VGyLtAF65cZ/9q71MOxnzTEWYtSDMCrO+JLHXnWjgJm2y4vYAnEA5
NzVRltEYh+cAZ1MKkgxzWHf3Df+jsYmjcYwgW43cT6/7KIduz1YjM9uQg+aBBrF0jJNA8viufzXu
blx9DV8gwZ9ezmUqpVLE4BQBRtkIGJsdAm2Yd3GYUSGc878+UCYaAHFVNjOF0TjsAEmfm+5rkG/0
S6bU4PsRGL08IWqJ6ai6BAloIEl/Ny4ySO5VHCbGrMiPldW44+/VOvkoDZ69lp5TlWT9NoORiWgo
JhSGv7fLf1TZClb1XeYIoXVhXkWWVUJA2aNLFEGVNwWWEEt35HkU2i0pcF318dendbce8vu6ODg8
YvGiD6wq6m6J6iIkYOh6obEGa9STLvmzut+8LcGtCUZ6mCkav3Jq5Aivp3quV+Sde80raaAGvh49
7nwaFBRI/ZUYrDvigTCB6Y4ZAOX7c8N+aAFHBpWAZl1hBY8Mi5n8S/ZFBM0601zT+5mjmA4Zlrwe
hxO5YwFYn6n+b4k5u8DEiMR1U27NyoGau9MVSIy0CqDAd8rsLrx+tFIAS+o4rlQX5ESGrAyEXQ2w
QiEZSoQLlq7MPEkZjIJbM4fg2AGo/f/vUFQJYzfjDaMFsqIo1gUrmvyzKP29LGVudrF2ij1fc8X2
xvHcGnyR95MP3Rp97sLKPi2AafOUSjsHpPA884aApglFSs4Q5zm66ShFTRHzZECUexn0KJ5nu8Cp
OLmkDW9TJUsQ4JbsKKUMActeYYvngNGpXdS3md0FPRxZhFe9b5DnanG/TIkEqGtN9k0Pk/bwmQ3c
0XbgpoILIK2VD2zOTYvLs5tSwTf+xXanTzHSgOEwxZ3ucg5844kN7xyEgEFu9ZGSc17QqT2++EZk
fG6gR4be0EgvpZlqwoFMPIiJCyC2MtD9F38AfbeLdjcdOZwhhws2e9ZAE3gNt9xEyi9sr2NS/p+A
PWt9rSyY/kLDKzt6FTwtpNxf3Uga7dhO/3lq0Nfwv38cP8z/SI3mFVX9bSQmXsiYa+6KtFp5l9pA
2GlIezakF/NHOD8nfSvPZRV7Hxqse51BBEv2mgS5Odh6k5YMiN0sSPCPHe2G/KCet+2lnZ8jPQZP
uaiTKJoLZaU8DDPkVaz1DA85FFBMuniptxgbEXInCpWA5zp6w5xM7Mn3bsxSqSCEGc8rb142smu0
LJ4sFaEwRb8Gpe2xhHSc/dInSExZq2oeLL6hICguPwwW2FO3HZjAVVpl2KTOEs4OJOOro3ZEjwIY
MLJulsAcnHvm44tKCQWBbNSRTJeSuJ/YRx/0O0X9ZuaSbpc8LJSg7QbCU/OJWmVVE1ntYisqLfSf
nzuXhaj3aWY+m9wO5/ifcQHeO8T+7Tr1NRiTY8E/L8B9FpibEIOoA0/+MAgK2rNXsWx8CMA53184
nHPcHw0JmWEtUxmEWKeeeFbXoqj3LhWPaXFzJLCo2mhcSVWH18XDr9geUjg6xMEytXlOJGI8gNY0
vO2C3/GN5bU/urvtAG5vOXeF23MGztp86s2a6J+MkOitqa8PLrIPqG5SddddJsAzYCtSKCFYyLer
Jzp/OgHPfs/jBpWw2D86eZG3P+9Jg538wDrWftNnuCXtUV30pyaQi9OUpa43Emk56eUOfN6amL0S
RYqF3mXnPemncLeQ96d6InFYSQJd1IK1ELghj7tDoa5WDgoQ61aFeVWQea22bqkzk8A5JEtLmHSc
u6jqBGBw9Gbd5YfV8+M8jz8p2y72ap9wIZiRozkk1Wv5Lnus58mSPwNKXgN9b7lJ2gg4O8xCFoS6
XHplJV2nwrrArUrzOV6/g3SQOVL3CONNUIy97SxvAnCHO9sOtNXNds9hNILL6/JKH863IkXoVknG
EDvQu7iJPRwQCHEMZCKZcxhWOaxGuQu8UHa+J4gfKg41AfptR5nTJwkIURHFRupipt2IJ3HyOAF2
isKbbAGTRJk7SuB1x9kpMtlXj6tE5qou6NnMdlRLX3Ggcf4l/4hTIVI+xHSkoF+suvervThV/Zy9
YCx0KcDcjLKthMI7AopMZLsTE1ljzrrrdaDByFNAggLiIPtkp+rkmg0f+/k9iEDpwYCj76MVF+mv
rLLt6XJVbr3HiUyZpiVmLmm8pG5Qhq/n7Dk6PZ90/uGYSoMPfie1sgBZAtKN/fAQ9eRQYXy/peNX
ibYaxQZPNQakjCJxKHbiIp8EZXCDcgzbfR1MlrG7tSPXKD/v3vTGSQ/yDZM+hIM182I3d+KKF5QD
tNOPy1Nl9rqrXf/e5HUFnJQXXMkRTogIfWWI+yKoZxv9C16jcx6s34jbghAzyFOMJivdwmTnEfeg
xh3W75YbPNtsdrvzThFR3zBLUGo/cNVlzHoqGGxUS0LjWsUXTyO60sj3dAzwpYRdWa52pmAPWYil
ry0ZQkBE+TRZmBRXOwnvosUW6ctIow9zua8+INtSLSQzSqZRsduThW8/g+WKBStPO1GQt6sYAhRg
DgBdfKWkyEQwlER62YqV1Va5RYSwMsQDOB258t0iwz57ieYq6KEuJXrcmQNxzOw7DDyRSW0GD/WD
0/5N4EaWBy7O5p/jbLO3oYXvn2v4dhGgI4XCqD6z9xm9lNY2qd5VxpzFxEDzxozRZda+1OB1pOIZ
X4gp32dDZZSZHaouysTyAGLBoyTZYY5peBva/rsHZKwpEwhRDwkrhQHImC7Ew+KrnOH+VzBOa0im
G+pt0PPBL4rN0Ypt9GUOxN0ni+AV4NABoAmaBgPOajhZN6aOMRw0+opKLrQxKT4t8IIYRkkWT4oo
cDAXP6dRZRtkjanjBajQtBER3m+PjGGkaqLWwJHSGxmU74CCQGxOUa5pfiwjRlO5wnwC/LFVZnUK
wdw1uh8yoXKcZUNJqffd7KqB61J8aW0RjhvRuR+BR3ciHPUDaXMw0yf0mDWRMlsqldYv9Zb2bdpC
vQ26zfDha481nx6/SPfpBO36rx6YhhFP3+d1LxjovLToItX5rj4xdkydMIPvIu+0fA1i3/Qa+79f
I8MOMGap8zeUowRjGq59RUlxIb6Ce6+U6QMpp6S99AayDT5TkCAV0zHzpqG6wyavfLqe4golwsGl
gMOfVHQh9Q6Li+pdTyMV1gLwHv5fXmlRaDGh9qvwcFTWhcUitRFuvQTLBT/MZUhYNEVM6aE+gnR+
EEwxiYkBORrXCx1ZtxrjTpUQljeZIDYgwoRLbdFWbBzegN0p/iUV2KGLzm1Hz9VRSr3YfK//sHp7
eqxsgCKm6gZAr3EwREcjDI9Rw6i08zpZdi5DAPIwQEiGZyAYcc6/c2vnnmdYBXgTChqvFKvya6d8
5WLSOCzesAhhohf8O2H8AtczgQ0QdM4KiQwCeFjoQMUc1IV+hQZX11iUIw6Fvh92JAV2cOqiY6aE
y6ViPdH52SUx3jMG2b8MslkdtsjCy9Fmd14m+cPmbj/P+//CyeznZjnTFhArb51fs2f0vKyj12DF
n3lXE39tXi0mkJ+5RRoW3UD1Zle4ITIU0urK2fhFZ7GAGoy0Jmuig7/iOBj2vjtgn81UQbww5/s1
D8XRxD43SpMnEGXj6Mw8Z58MqZtGWQO5lgpnx2Mx1UpTHA0tdFq+wcSx808wQxADGg5/cI1lku3h
PZ+J7AQLQvWhe3oy2+s1R+M+EyYMgv7/r/ukjj4mYCn+nz2OOtUrnW0XxcJ2yhQ1cH9A93uugQGh
DcFCbpGyJEufjEMT0YexexmhDx7mBRljRsNW0BSCgAaXAw7TIlubBKoOIXjkqvFRG4kuK+5rh5Jx
98NG1len7+hVYEKretixpJ6nnELFurl+cehRnslpzvZIXv0yaBJ8ksrtLlpepCqBHjSwgt+BNL9K
wVUQ5CG0fN1KFQ6BJtvF1hdyYeiNbixuC8gnYq5QRfcwEnLB/GxQOOUK7VH3MZI+Lsxbk84SNRTh
chXlfThzM8WJfGRGiKkqBBb5cevvyuSARqVAGuabr/88yhdEN8pDHy0uGKlWsNnVhoHnQempcXLT
KTy6dHAGAb5+/qU28GF9LSQbypJ2Txdnug6IflmRaw1JGBPb8hq47sFw2CcQyoARxAxcv08kKeyI
PWnbEkLa1MfUROi7sV0Boubyptq4e60QMPVMkii5gyqjROlULcvvM72WtPqghGPEEU04FesQ+2WB
cRlGYBkZqoyU+DQS9SYLUcs4jiebY4ti3oF8xeM2o0rMiBT5DEJscLMxXOnr7lcFDEuygvN7Gnor
KNhp1yO1bxVMMUkwKXxLlwEbCLF5ZvKPx7msa2SfsiB/w+b2ZfniFtC441vTBX5tD1ZOcYB5i1b7
uAYRKaIDrHYEQpeBRbcHZeWh9oH5xinL718F2vkhZbYgUNbx+Kc1EtAnShDgzzRb6F7hWWJ2AgIM
jiLYgNY6LGg6ReWk5lJm74EZzZOzNIg/jlkytNLxDY12OUmRfdm+zzjzQoSOuPgv5khsv1Vmyo/V
rzTtlCOG67S/GRo04Qjfduz+Xn6SKns6aN3DmJ50xBmWHJFWPECBiRHDAFCyc1bkVPrhioMZ0Qbv
6OYmb8BNTRDRnVl4m9G6cqlSsMbFq5ES7XPTlWC2OJLMzNZIIohJEL0c3oQ4Ic7/WgP19fD6rc3e
LPQrtVDhA2MXFW1LDU0mGF0AUKxzpxOcgAntizzemmLW7syNBRE0YwT8EVgZY+Bjj41iPlP6kaoF
D/aNnTbRNavsSST+wyC9WFWKLPFXYItsNQNmqIAQIQb5nPSnnTgUyb0tax6k1mVwHbfr5G7t4zeY
ZMsI6XQJzLYcMRz9UJI8/nT0eeyGR3xPdp8/H82T+SSpnROecqKq6SsvaPqaJuUuqaDnLbx01fRk
OPSvXh0Z+c5I6x6IMKDo8bS4F26Y9v2fqLBiTqCkcToz9n0DmuH+G9g4Z/9RpabfPFUViTmJQLRu
8Pbc8nlOtsdnMi1+HYBdzwjZvqC+cDmHm9W+tWhPekcgYv/nYRnCJysxBaF3Oi4+8N0n/NWRBxVl
kaQxgyd3O/DRfof5F8CH8tFkiyh3bcJM9H7Ne7MgF6SLgLt+VdPSGleqFNC2Uae7+w5fLQLIMqAj
qvAsHsikIgISzNovPQonS7CAqHd9m+pLn4BGFjSs4JEnW8BU7bA45AvPM4vS4CUmNFwW7yI5Gybe
aj6zSbRGFNGZNn/SseXYbaQc8QGbQDXRP7allVLlqQhkH1eigy4AvcGmZVhcajef2DD0mI9grc1Q
mwI8MzMIcaukbYwu35jSw0g1RTMKz/gDeo2vQxjCeBSFXu1p92gDaTbnj2ewqR1PIwHtumOYu8oK
0b6kygoSVpGGiuEfRF6aOrcGHNK5cIAGMWOGx/V8FYAIl8LUWkmBN1DZoGp72y/Tdi90VIPJtEoz
rfh+OyX6dygnQFL/rivgHVLjj+CCF36tWo/1xaxkxpmQTOiviNjhMuGEO8YNVC89Odp/u7VU9web
tr7Ph6QwjO1DlziHvZdsMuqNtg2J4dR1RJPTqWyPLeaJNRU5ivOqkCFSbgvfWhQb7L4QAy2tw2m3
/fkzq1b/LtPiA96dgpkkuThmd9+LQGtdlNkkRh53yXpPpc4xHtlyKuVgbGuo1pecumiCH1duqTtH
9arr26cxDWFVUncv9Bz2l1CmkyHfqQeT83snpWdRNW/xA+DfgNQ5/HPZtFcI9ji34ywu1tAWRjRh
EOSe/AY/MsnX9dCqdyffsNn2CCkUiXLXmzBF8LgNBPOcLqx3SEs1fl7ZEO9Cl1tGCEALv9VTEf1M
3CWqi0moLr7gH1wrqMjEzBKJve5wlMDMlQlGINL6fSl/eyjJx2RJYdLI7s7/FHvE1q48PjC394Tr
Cw0hEliXrHkJnsA8yCeLx+avzF6XdfTQeD8cKLnjMZJIyGOhSlEcx2bHIqcchwhl6hFaha2+ybeu
hQjrXLC55yhLJwNtb2XmAVfi+xTYDfrOkSw+M1oDmOl5g4HqE5e5CmsJiT9EpCYqZz+ag2c5r101
sneuvEtijiEz7jrypGg8UX5QT2OgTzgYA98e6TNWNKLGdCS2RpySg+bPEP9YHo210dHwJg5EJG/x
8rb6gfKlhpZEKQ0AhkTfubLPwIX4bCy8+x+l0rKLOt7TqOu+evH6H3lxzau82sNYQRHAVaFFYgNP
osKovIDjg5aOr3O/5meTbv+wx6lgw5H61IVHfPYvoeZRT8mFF0geS4npyGcXSKhDBddpYU5y9n7G
jsJS9Isx62zKUv6c8SCtbO0jEnTgoQB8Dbx9DmuvMtOz8+UGkQiJ767EFL+4AN4KHsDk0sdKnF9I
pVUSPdluCWL1sF6aI+z8oZ5SnV86F4UWLs8E02VKKyMNynwaDgg/nXJAkkfO2BJa0mgmeQyoosoX
wwGK1B1hbLHLfPMqE0VhUs7UpbDWDXC82XlgJYv71RLoXqbhX2hZFBk+iiNoLc4OelpOIRnv7Yde
dVEgWF/zG7WNYrp7zqMAWTTO6FPm5K+aYUPxSg+WJBhKZKqBtWNIdRd4E/TnXrbtV6toZfktUkvh
hoJIUg56bHgUzU9uW1Ilp69Edbx7csTrJvlAammZnDYjVJ7U9bvn9YUV3QsA39Rj1rXcAA2IS+Us
ZVmaHqLB6z/htRCSVqe0y2uK85qKMagN/3vE5qI59hCxSLm0sPV+00PdD+r+wFlQbcIXYKSrdfhb
UGepROMvqu4F+YqDGeDlgK0tXSCkHo/Jqydud+NRoAmno7Mt1Y4RgYQP+6/kgS5/hVxPT9v4JXRy
PF2vHCUhlXR11Lijyj2L9n5QGzaSz7jlGydXV+RDWKvmdwbVZ8r6CIOG7/Rn/ngl2lGN8cwfjAAB
ePFEF3QD3qLZ0K1kjCA1Pe7DHJaRIlegYqIujmPy5Y+qQ5Cg8CjfamjBCn/DIjKEomRXCRGqPDC9
ERxFhGKter0bHA1/T+caj+3JbttnLIUFdkHKr7MbzATGh3AfIe2CM/KFact0OtABR4s0lvDSv8mp
PMHw3LuDqMcRFER93EE1MgI5Om8TMCI66VSc5aPMwYpNTGnpr5yBQO7K2MuaeoPO0KhQLaivdKij
bSknTLWqSfkBL5txZgouALuaZc/AjvxkprBv37XjWRAcwSna9oMTZCsOx8AK0u34+Y3Z5sAHX4Ge
x8RmpWi+0BHkDJ5kOHiJfR0JDDzwCIHucIt+PB4PdS4jU+Fn8UbHci5Osw2+AkwFKGCOYxSr7duR
4E2KkMIThySx2VUWYdxN7QzGLh9r2FHWDbPAZTgm8SF41YmwGOo1i8DMQatVOEEaO673igU8fMe/
fNCFBzrlhaf1OhuCL2RBV1bJmdiaTuoGns1HL6xz7gKCVZ6BlI4TlNOP8AVrFQGrNg0+9nCpSMwS
dedyUXDy/YpbqdJQKLCMpTzmP83O9awFnM6ypiHUHmp7EqBPSyMLo+OJ4hADBLswT7TuBFRVGerZ
Gr+6MWdGg543AB8UeJbozyMg21qZc1WeZw1/WJ1P6n4PtL/z9HMGwynpMW2OU8xLIZ64oX8LXZ6m
z7+MDgJ92bODLws2B/l01k8d9CUGxUuSz30S7X3JtxyCpmgUjKAf9FgN1mRdtenlJf2vOFlYq12s
CazWVAhsQc94UaVOizFa+HYq4FEtHQJIvZTZdGK6+jvXjjqGCUdO4+vvXaofoIhF5uEFCIrqo4+C
Jyk94SuNT+Q21zVsxTUALcl4iQkv3Uj7Pywdv6Ft2NUeSf5gWUbXpbLSL+I5tUbb8JMMgrpWDtmF
1s46jcTSkQasyPvgHFhofjqpIfkZnn7RiOrK9A75bj8Nyx29JPARHqIvEkoD9XxlQqBOjE66iVn+
X9SpCLSb2+eG4TtRjNGGJaxo/LwvCxzeJ6KfxdvFrOt8bWyEwnCmjV7+YfZiIYeRXtbf1eztHWAP
7vRrdD76enFpxiBC6wWdfxPqLv1x+DyHctcB0dGw/jHIIawC5cPfdB9ukiOd13dM0F2OUgteItXi
qGHB28vf0r4z/JRWn3QxFRKtUwR4P/5UmwC9ToJGFFes8X+/2nUZ5bEChmvEpeFiQcIZAlhIMxxl
9/n6A1w0BqkXRSVdUYbBKu4oVMmPGzskAiDqnqbtUD2tGTLhf8cClbfvbau/G7X+H1npVvkni8sN
mtck8ap8yLNP22QorbOgoQIXtVDdrMU0eMF5SDF8ZgyTaqfX+kuVOgsM08OUQTl8UKXO9F1GRYIw
FWGF1m+SWyjGqHqZhtxYp/T26R2JLaHAsZK1X+BYL+iX+U2bN/V6JjOyeJVdCtKOlFgSP79/3AEh
emrvrUMHIvkI6vcepblifcZE8JvqdS4SgUxSoEBgZS0tcLA7lDnG9Z6vv16wTqqmXuiUhtxHhYKk
o0l3SBhwB16EZD6rglVEoRT1Jrn2rstNPK8dzOV2hOMr3nq+On/gDopUuFomvi3IbKw8JEF/YuV3
2QPNGwzbUq7sGtKF++NPTw4AHh8lxCHdJ/jy2HYBHWNg2L2nJSMPscsCGbtoK2GZL+90SS52uxLV
NNR0uLZlqVISEoMjTin0l4BTqRU8OXN5w2LqAK+Ypw9NGJjYBwlboioQQ8T4L5dXM6zFaSV1b8qF
OQ06lJARuwPvxbu+2nWvrXcKM1yy9+J2iQQkvrFTDs/1Za4MI6mKwEUQXBDfKmtjtkeqo2y36St3
pPAMZZkVIJxp8TfgivM1aZcGWReZHaCvaAgkXAwzkefYRjVs/dHcR/3mHHTwToBo+XypZYmgyIK8
QmGZ6mJvlWoHrIMtQrct9c+1y2RbwL7O+38Qveq1dLy21AadaO1xF/JDIJD3H9/A3HPNHj+AoZ+u
xc8NnwZcIjV1JefScQESj9Fe7OnHiitSsV5GgyHjwZDcFmYLhuKMRiTZ+aEGt7DvHZQUhJ3LEh9N
NYNvIl6reNofU67quJGl4tV70ocS/jbjCuJn70LlekrUyjOWunKqw4iMpYS8W4DcN6Cxw0mx7vH/
4D7mzA3S9C4xAlKL1cVRKzqarR9Kaq3KepYlopClfOabwuwpvjv2+MkpeSFQUXkkGJ1dQrYxVkT1
mtYmrWEVAv86IkxE4wE6BUJRmzvfRD2Vr9btGIptS9gWl7grA81sSZBnQrYiiypmrz8M+RJqY4xC
tJNtefY6+jLEotnuQm/oiXaifxP+UOEUSqSTc192jP2yRPRx6KEl1+IXqPPZ2bWIk+063CqaleJK
cNupgQ8C4B0OllTzYWw0Ldq0T1D3pxJRFyG511txCXoDe+wG7L5J6ThrKMuFNRM44xusXeFfX/Tp
C4iq7ermgE7v5O8doYNP3VGGC/TEI//T3MhKt1pQGNWB1x4fuxuv2INbrknohH8mH4rVNnd3gPFH
yUab/CeFOAeR3W/PegBVT/D+DZSqsfBUOvsNslTHCh0LSvXZs0Qc59gof3EVA2NVVmCETCVARxaY
2NKVQCB07/UOLMNxWNDkKGo1GdpD6CIJKVDbyeQRBTWzSFrwhHZJCD1j5TxyhtJSI0VmtpcrM5Hi
VTSJsssZKflALKAsZNEfwoa7qy/Y4eLxPFUti5mhk4p9nIwgI+Q5VwIytMv61SuCl5vxjzIj6Zwi
/RWnwVLC6Q+aBnNyt9llysaBImHdox1xwQQtPxZWwb7o/oQaJUU5fQv/vNhBvRY/QPsv34luWLDg
ZKZr4afwY/2KNkEqUYRW01OMHeBChjpcrlLFkGLOXI1SBlDCbkquPDb80TXTPk7hepkzn0EWJlSF
HgWcJxkbrkmumhZErad81Gdi049OTUi2CpZhyzUqfa5ZirsUKAiIwkl6qFw7KQOU4Xu+b/q0Q0/W
MuPTtxCY8VIymeInVt9yiJE+k6A9OMZmIEstzSnbVwmqmZd2ZNit7F3L9I5PL+ivh2UCCytKbNRp
ej+2ZHxIdNw2rA6qOD3oeIRG/qtxv4cKOEXgsoVBfznnAhNddX/2jS8mNUIJzl21alpE/hk5hdHs
Nwb1c0Npkf6yFyiVDkp45BEFPdSgP+cbMV7dHroP2mDdmKzkUdryOc9FAxu/oybrQCnhJxsavBsE
72t1F4FlO2WELQK3zXknEv7CT/8sLji1eIjYiymHXmpclvTMAPjcIYPdeoxT+4Gd5YyO2gEmQ1KM
RuvVanAF6s3J8VJ3gl9qUjMXSe1a6+DYZ40kwm5oaVx2eDayMg8lTRNulaJAb607egOsk1N9pl/z
Uram9SSXm4hBhWsuvCvrlN4oFRZkQYxH1p6a3Dis58xFtEuN6QkM+R6VQouyqUYoj3URqQB4Kldk
ztEZ/pQ20RMIgoF0L02jvgylPxj6W3DJg3CP9i1IZGVnhPmFjVynPG8og3Nre8Q+SFsVPIP2NaTr
SQTDXNrI80wV5wx96gbWWV4bQG2//SScjLgwca3/StQbkjLkHhjCrqe+sNbjDlzkFpDh2lhSMSJp
OWkTIQZNZaI2afy6qrGgm5DC9MzeHcQA8cFL6SxrITqAcx9qKTFv664g4mxwiuQdZOaqBIBSq6Je
HuA4jUd3pNrTHHfZUG2CD7x7MKEqtu+S6jLEJY0UsL+oxYbp7C80RfpVfa9crPWXX9EsKZdQIj0g
xetrpRIGbu+HKyDXQ9ahFKnuluSbqkikC8X5H8IkTw4gy55lYQVXyKmdNb2iGcxazsLz+gtCRxKd
14Yldyd+SJl/F8ApgcK9SjvHI/c7TuamLJltVRS9ngTyG/b5TYbWuAvIY0K8TVdG5LRHRX1NSQj3
DjCIhuCPrZuBiAXTKpuv7KJ4aRnzLRHsw3cP93Lnkmk1xQeguUdMmVJtyzC0UKorxwZFSPGf67A8
r3iKD4k7yy93nmQ+jT/499/gcgfu2PfUOdgXvDtssy5gjNrb8iTTaArULnad1LEqCEwK2SuC0iol
4Rfxkzp5dPVjMRYFtPr3u/XHKKj4RhaDtO8A3huGmIvRcl6XcD2AAUUPlhy/cv1KAEDXjwJOEZjW
v5K+fH+16gXq76G+t8KyWmvcND7Zar0oge7Tmr7lN7V7AddxqI+RiwPSi4BNzBqN7PfGhuu6n8JG
WdtR5vBsGzCgT4uarEO5KkFMPKqj5z8gs/8YpfCdW/uPLrJCGq4rK6gjjI+/v4nd0zDZj5201fNS
eYZNQwitGbeFyi5+wCsdexEkfTaPTsB3qcYXq4jK+TShjVxYpSRY2OeHu2B2TcvfxAIjC2i56/99
geHAw/90t0c4+/pnJ6jQpDB+XPxiMrt8WUL38oeK78PjCsXqO91lCfllJcXAftosGqbaoxw01kgd
aMDrPItUS4MSjd3bS3yJl88Q1kJ0ATRcxAmNSbBl5gkb3mtwLzwSwwDR1PnjJIpunhf0inx/E7we
kbOD3cqiEx+Zw52ZDLbTcIUbyMNPAdwZEn9G+/TB3VI5Cgpzt1w+4jlplK1YBuwG88okFuPtf1A5
hwUgc/1bV68k/fSc9++X8Ln9TI22+EUFK57yDW+x5J7dStvzjFBhfvvTHww5gIc+KTDg7F82T9Gm
JUvMTvRpf+IneTzNlD4LJHo7GlWmbhc9zuJXvlVtXeMmmjogiv19dXc+Gv8iA6IcrKzmT9+KXq+s
9Zic5hFcRqvQJiPQBQT9TsZ9wi3NVtjcyeTyaikSzk3ThoF19ekkSXPBXm9e4L49NnV3Vq5JQAhT
PyaIqBu/yQSahgJP1l6JEfd3aunC0t2SCnqy0yGvn2Nb0ROrB+EAGxeDw0l3JNaQhrs2xuSaP4Yl
9CPrsylfZuQPN3Svv74evvXx3f4xO9Ib9L4vnQQlGXf6P4c/sxu19QFMQAL6NYqkq/XpDWkIwkBK
Lup0ij0PdHpQRxzlHyf7XKheiKBjPhzn3AwaHXlaiW/Hiy2wDCclqk+ccMGx/Npkg45RjtLm1Naz
eL0bqDSRjravPasXeDzQgHNbQWSSpM5qfwTy6FPL5xsnwUj1UtUUr4Wme4KC+w/q4qr5Mlk/aaBi
Jc5K/gcKKSYZEndx8xzouiLbGB+HGjpXBwFAxWCqXplv1nuQJ/cj2jOAEMn7BYEwj/AWAubpX3mv
6S/THKA+2vDGVt12E53Z6V0RgOoLf/9VYg8Gt9o2C21bui+VBJdgAFff3w/bqPYAJ/mg2rO5bxHU
qInNDNGaHb9a301+yhvp5xgiU36ryoRxYBHS+AxheqKzuk5sHe1fD5wTY6J9ylGgwECnrB43b958
0hBAH8IWp3j1v/nOpP3BO0MfYlgbCjAZxVhPURSdih9gzaNpJMctBBR9iitJBGMlMTL6mDqYdH3M
YVN4hMe3tfZ8GZXsf0wXdrzGjgSQDfb7a5Sx5CUaZa+1fgXenrg6dy8CRoyrOZrJqqMkYyLeBthu
arOcpB/Fxc7vtyfwzxcTDYaMMoQK8AQNCkTgEiImuO3WIyL2edVEc68DujdJajcB+Wv0wKeHcHrp
kkURHkrdQKXcqORuVL/aK5xbX5eFUMvHyzJz103EtrvpNUspMwbcX8+9+iGH+xmoy/ay7grVd3dy
JCWyznaohjtzo4FDBKGnBh5WyFPCag+TzC+DMZB85W/DpgFEBas+HCBwOaGGId23EHdC4KmxXzL5
c6YKZIfsf6GxVbMMpSobH+z1Z0MhAGapf3ofxqxLnZ+ia+BYn3/WdCpeGsUSNFNHzSFkWdzQMxtP
tifRfa5/cq6mQXfXbpjwMP4oraB5sCbaMqdijFJjbZy2BtGmBBl5FelhJe/rvGA9E5ci6YCJR/Q1
43BulNvRC5MDigIp1VzIYHHGrjN/8p5bavWjFB9+T+D8gG8wYRqwZwaZMFQcKAUjhXwTQ/gLJ9y+
9gHkNoYSQEYl+a7nz5EAXXnnlgG0VaiD35WdrSMW7Yb1T5nHrQb9SuR2o1rk43pxALtbSOpuMCyo
G9OqeboRG9d/z7TTDKzjNjkGCeXPIwo63ogS6sgRnc+gtHT+GgpFsFynSC5Z8ROlHg8nRZ6UUIah
1zKSrJzP5tk4d+ztW3BOBUaOD0JcqAVCVeN1XmcqLCZ2a4gLebnC48hJnDJG38iaqazuO90fAC3m
55UKvH/Yje2KyAPxa8L0IooUwWIfaAOD61p7RkReZlwiKhAUXbIW6TdInMHdyYTBbqSoYD0KNnCQ
A6hEL1XN5Qrb/IDhoi6m5pZ6sNkeql0Foyt0ZvGVY3CZj8QGtybgW58tCQ45MUpQ0D7mjMif02Ty
L3XQN4GZQ/+uyFew8l9M3Ye5j/y65P4DoKbYgqj4fjD2J7g3UQxGC/ungrpGmVqEXFOXnM+JHcNG
yvDE6N7lw69smUYu1QpiAvHYpnmYofin+TvoL2/EoyjLzLJM+2PQOv4Mf6GANiFu8qTd22vTyLwz
WmyWNZA3V+FTQdB14Dk01uXZw3fTo3QNtrP0Y3KVNpfMsLO6np2eQ1PZvI/mdEPBJkpL5xFIbt5F
xYDok2SD5SeCsw+sPgyY4ixSj8qm/YhTZ+b6cDdzIAmlHNtgjO4GhNlVSBCxrPJBRSjClD0gsoy9
Gt+6/5VvLslV7PdiyZ3nOxkgjeaiDK2xdILwcYzQNEkRzx0Z91BeRQASytKwJ6AJNTkCjvq/lDvt
7TzLNIkyqM3ECQ25sQ/DWSTh80HhgwohmLQkY/SuMbfxN+MUhulZBc0LGexW0X9tRsk+J4OjG8GB
t3dNpt1Mmq9teOhaH/HmR4qOJp3tJs/8AwS2pa8LkFuLHomBpTDKvB8jvfNfx1+qIpoqRPbMs4rC
/SVyCoIwuePCtJUcnbsIbjDmDsXxajUwNiEKoBWyZexmay4dIDtgvZz/hvlq2XYuw+jVJEJzAE0w
ACv8ezEoali2k/J2MJWnZfxzTx2x0jZaCPUxyyVU4b1C0kR3uKCnSD8WuxYWeuGmiOtN5e131n0f
QK2pEmGU9TPzDbdPpdzMnoOltm+qai/zKuOFZtZX6yn8IP+y3qm6GgzQPUCsi3SSe+uYzV1vc3af
WtjDsc5F5ZR+Al+jQkUID21vn19hUdMculNF7NFxsqMvaqqBFZo6iST8ElC/Br3h1Ci8x9XcxvAC
JvInVEcTznep3n5cWIsrB9l9b5Cg6f9LyzHJzxJ3KRz+iNuuwZe3KQ6f2JqehEyxELOtn4CnnbQd
GprSjfx3DI0ZS1h5x/c3bB8pB5+UyE6jC771/VxEccOoK8oc0Veb6dd1t4iWxz4naGxA281NeXNw
zVxBT5s5tw1wq5FQVYQMvFyOl57NK7U4+L6AzMS3G6ei94LjGheFlKTFDT1uNXmipPN5NEsq10Rq
7gDpPADItp87eCYnjNwfAuNSBWtp6XvI7sVuVPVOitXXN0YfszBpuhVeawxNJhI8ZphwkgKdoVRB
NjyGK02nSqdk9QJnDy6sUTdVlcW897I4jSpEJeFjCmltsR6WmwWMxW2m9o0sT87Ea9aaZga/s83f
pW/NLF9Mgix1SbDI6H2Mcx6SDuCXvHnKGCZOwbk48bZ+3vSnhm/6gEq+R77RmaOaEb7gecGI8reL
t+MSuo89pYasKAe+A2va3ESte8JvgdfF/y0Wno/EwI9lWVI8CFlW+YyHjOd/95D+DGLUHbIusq9B
bYmgycoULzLkRWpZZn5WZ+RDYpxsTphGHGyy61rfvi3GPblQ19EQ/nr9XdHFVTW/OaqM2r9zGVXB
sPholZbQnznh9uA5LaDu7yzsJpQHYr7AGzgb5oxogGBe3Hr/LNvZ1uCDsuFRU9LQln956fY2vwfR
ckjxD3kxuexIgTBQ2rK/K1zlAJOAOJjo+UpmhVBakNKpV17b/PaMsoo9An9fPFSjbm0RsN4oqU0g
xe1kRMCjPfsMMVSLWhdfLNQ9h4y/jWf0drsZ5rTtLJBb5/y8EYzXD/WjmJ4qvNLpfrgMY1GHFMAx
HmSH7ikMdO45BKAyCQgNBKn6rcBReDa/V3CVKBWd9f2P4SiQZg8kGs0apPlY1NmOQx6bJ8Gf2RmG
v1SsxZkj5ok0VruMf8my0ApdZD9POAXL6zYpDSshxgON/0oA5M/yQuaMdmfl+LesVsFQlPbd4S5x
cVlqOGTRUL34uafaMqcjYVcJbxIN6regYYzktqcqO62NTJsfI1Xp31QBiHBHgE5v0bB4pRoGSgbv
g7buxM0W6tADBvemtbktrzpDRkmwkMCRHwLwoitEiQFdTRS7QmFLodtuceeoJiAm5UTcQZ6wvUSG
ACnCwaCFipRwh4aOhhAxYdnEmzuzpX2FnwxMgdgsYh1rjMR4TwI4lEVlrWaK2jfR27XMZIkF74zI
bt9gKUN9KkhAyd5akAG0jqKGRfkns3tiOddVuDXgHTs4BFOqzHXvK34kmF6mA68ok8ugSmd5uzay
wcw/q5CWX+79FhmrkDKm8WVixL9RhQSGzWokqdl2e/BQ+FoXMictVWvR/pFDorMVJTG5gtuLE5L8
OBokWj+0uDOuJYsim67Eh5tNXVAN08NQu9tuCdVHJA0vLDzuqzudmIbmxwStEE2dNqB1D41rmJjB
e5Pi7aylb63o+TAFYLDB9po6FKBBrRTSQmPohZDmW/2uIR8iJWCV60PBGsHrqV2HnAwE9TNL0f8V
h3Jt7edDowoKaF3nvBQCIjDqhYtASwqn6QlFklszQKeYu16X+FR4P96Jgchdy/7DLgAkoGisr993
AXgF8iMxiNcVUx3o4pMaclsK6xp6Cq4cZx2q+r6V1tyQ62LpdOd4LP/CKnpgki4awDjYBtyl4T1d
tUyjvmHUq0Csa4TsWETP6ub9dEHxxUHJVl+mgpPsb8fZSZe2d0b8ZWEb4lBKOllu9eeqRa/C+7I/
Up8MUtu2+BRO7GVuUjKSrGVpV86aHqlUWOHhBOLJOnP/Fz/qEAe3CbJtRItk7s6HgP26+/tLZbkL
xFtMFWIflInOVwiOd/jKT5bvGVUd3eQ/VeSGepMAN8giau/7DtvzvwbzytANd0XKqJgW1MT7yotD
DA4bwGSdQfsed/vMvUZAQEFLVg4p9X73kD4nWLtytpTOC1TjW1QBnmvqJJg630AGg+kVLElKZNvI
VgAL7gZtbAeMZdNKcP3ZaVea3+RQOTuQuBwGYrThM2+i4eZV3iF/fjkXG+nE/PDCiyy2BmmjO4TK
WP5W9mlf0k3MaclJVRg9RTK7I8Gsy7XPXSW7XkdwMcFG8KxZkFl2NY+dKKhofurABjbqfb7bB7e2
i4urjxWOXTHcX52KinrZoV5gX4ApN+/2NWEtcv48rff4nXngZS3vCBbBQiMlXMf7cRLI5EUBC6c9
jS9Y/jl5Ik2v3dwNUFcIFy7sjkF73JO+T2iS/Zwbd4Kag8SHi3EihMwoKfJvwFnWFtniQaWb7W3b
p7duJZLQX/Tt2QQcjrYhj8aBNypLL7zHzP8IxXrOW460ZS3XZ09YWaV0QqhwN4n4Zuu303JEOSlq
sOoBH3HqCNGxS0lZHvHdkYfoR4wKA3YwZi4fkbVMVIIqCwPqD0Z60K/6bWMMA/g6/eCM5mcC9LKD
dsA0HIpBBjp+ZdFFPqc1XPJKo/B/lb0EXTs3JwHo/e+xGEet2V9bayotN4ibrl0UFa5sWaqjWRzx
Nwi6vZDQ2WfXhjQ3in7rIhAqiyBiwiDg01P49yXdPSY/k47w3np/v35T+nMwABeKLKX7SE9oeoms
6oz+yEQhQVfuMlEreX6x3HYUGEmGstRh336i4I1l4qT7/O2PtGfA3Y6qCnBTP2qZbCRU+mWttyav
NkuK+2qhrtbB/seOx7PcaOJ4h5zLLDWiET9JwFG2QXLsQ/UMhywofCsHM1dS36BwYNGPDqt98eRg
sXYGxZU5L2oonL0mIOgBJcqzGCC5oYB14cAVYSysFSK7QsAX4jeBABIewLQOBbiwBtYqKSmJWCKJ
ZgnqQHSikYJxKoAU+ZKviF2UJpjK/dFCjdudkXYr9ay06Kzkcygj6NmKParazWQOT4589dRvkBYH
cPXnZaUedd5NnLx18SGKZL9rz+pGmllBRRUa++NHmi0QmrGtMkrudAVBerq5Si2Nv7Ix2Vou+Adc
pCHeEeIPf73QXwSytMfZ8C7sqihCxQ2u3NsxyARVZgcGq5kXGS9jDaPxMKCRKy2fYxWKgaoh0xIm
vIJxEFKYwLyv5rLqS/pFUOhsoX43uIXvnvsnz6Lx5QSnncdyRM/B1E1OP+japndzdCANXzG4xdHe
ImyoV/vKRZ58eXDm2xfv/buq3K36lbNjuDQ4r9T2q7mSRHlz8iouy3ai97QJkXYC8DIFKp51OWeM
WKOjnUzonEoSXqQ7PkjJZzt1cawlYWqLb5pNGJ3AzT2s2qup56NP/ChKmPMwe0UzOVITiB6PP0OP
PEBBobtleNlOc+6hYyiGJlE6JJI4N1lVdJoVBRkO+ECAspmeEEXA61fH4TDnOfe2Move2jzUEM3t
MJjeXkVP/RDMStxXGN6nHQWAeyJ1JAKchyCeZNNlJs74YLqmAX0RhqpZHJl8N6wPGGo8dftH8axm
H9AZ99/VBlnXvvsvSeShIpddqMtEru8iTn8AQTCcC6eyL+Cbm2IzjL+h2qV7iPtQlVSgXwIXO4le
z+qbujr654xGQpTuYictP3xd2bR0BG6ghrRASt3/SMmdD+uBASwFE3DV1o8Xup8WNko18qJ8roEr
O0DFFebMFycevzMPaGkivs/FKpIdpt/cD1ytGzE5CQvJKfGFSNvwnJ61Ullktc/CwPE9cBd8vV2R
xxysdixf1cJjjzXhLs3qoQkYspgQ1FWXY1q4t34xCSEt5vzpGB4LIyfFwuKMmK3QZPTvdGTaWYbm
gsQTpUWUmZXWyDcNMFJPdHUx6bPFlqrn0wD0MkBNeGxdfZB8S/6Y2p8Tf5pY5nW7uUtj2m/yGf4y
cty1YwkwyEU42LGo5zrZbygSG42PKufw2+EhKhla/Ez8FxNM3PbgVAc4/CI3ay4Eqi/dUGzFDzXU
u8hSsOhDJnlSAFofikbegiJbeb9fa6qfBtNvXmr1I/Hw1EVuJPRNPqPSr76UlusA4oceBUwcnKis
OnKfo+PwTQR1bXBmrju3fr4tvREYdpRujfL6xFeB3e7wR35DQClECphnMGe23y6m+cUDcJOJ7nP8
p4H24OA8AxrTerFYE4K61OXNRCaO3rWBhLjlctyN+GPwoE12nMNPs/4QX1panhMzP3UxCQet09K+
gDL/M7apxztrdTdDuelbqaQ/RHEG1ghEDek/0LA+PBQLfc23Pe8hZnc2DwzvqiQN8I+GVmIXXpLA
cjkyWBRMuaNmm+k6mo6fXI1bCAoi4bddq5VCuphm1+jxHgWJwdoYlUGguIlk+NXA+zhP3RK6228O
/t/p7Dhs6iwzowuSYU02qLHCQnkTijUi6Hyn+gw07f7XoZjP6B2eJYMCs/xPAgq9BLjddbobyez9
pp+dCDW7GrdCEqnTYau59ErSTNRO9pcvEE64qrgi90jTPg9OM3pOZT3konhlG/e8zRa9yuwJInS9
F/wXnC9/63EpeJ2vBQin7UIos1zHCcCqTFbdfxU8LX0ECx3R5Ga1x1KhkrGenDv1N6Vd501h0mkg
m8VOn2qDKuitAGNyLxHdD1Tpk9VMjtVXECn1t+f8120vFzFmlSzCzmxnVAdPr+RSaUDKZDnp6Twv
Pf67YeRcMBXIwLB+Fww+HNxvPTSl3ENEyPbLPbiglaGfz646RcaOKfSVGSTMGUOp2PRh77YQHiTd
1XE8xaX7V45ZIexFNCgb/YFWIfL6Ho7TvsGRfQaI/Xqig/ECaNvQhN9jeLMzc6PsWSF1tzhb9A+Y
PleN+GW84unFV5+qSjzkRzkjSKHJt9aMrgKupRKIuRuyq/Io+xXi0NmTVuA8Xb+4UaCtqWQo1Lpc
+ThqUTVhQVnnGDoTwxtVkidxwRiHr6pL/L9CYYVPj97dSQrmsoLAq5tKQmOxl+mqnkxcDOHrp5dH
bo99+terrtlFH+n3WoY+9Y2sqakmmzStkzNPkK2rhv32RqxU4D4tIBUJXPgiNZJPEhFmHOAelsa9
CcVyzTiMO6Na0xhm7FXSN2htQS3yTbo3/ic/FVDo8GBJaJ1WHYf1ABARKXYSMUiIl6bEM1Bs49Kn
ruxLRG5H2nVwKTqSPwGJPaXkU4msuHtNexHP0wfWGc2TLLzLayvPWhLEpC1293NYJ7asI9/z+h5s
l8Y9D91vUGzXPI7PacjIUctH53jWDWXK1Y0bupp40II666E2NMNVz1UmDjxFxTreOCbKTiZRHrvH
mbm35L3W0Zjw6AjM9dBPAWvqWrTOE3jXQcuX7f35BqzaMBeYJI9AA9vDGvdiFMOYgV740TXgIHIy
THes2yyIIgSqtNyP5gRvk8gVgo06k3YhujQe8TizeTvtdMw1HZAA6zEZ6uzLl4pWea9sU4UKyaCh
uu2MojWeee2IgYrtE8k/aza6RIs4i7HzshoV3mgEtnW49Ek1DRhegU2Bl+joSW09p1AD6EpVP4/4
RFtsq1+RY24qAxNsOiX5uB78gj9tjDr79NoGaPeAjYXqqS/2Fs5kVE9mxF0A+N62p1IIx37Q1K4R
MOi4pw/FgagPu6kUgqESZU6iWJdXK7kTElOapCixwbqAkc3o4RxThu//yd5FZkTRRtsFeTtQwiwt
yuDbHCe/swfkd5soAn5s/cAC/s6+nfLGEKkrdvZ2oP0rqMpJL6PwceIJ+MNOkK4wV0K5Yy+FF2jI
NL9RBTK70NFLrGhXyUC/Ekc1id5uwQDT0aoidnsxnjZwERHuj6spFWpEZ5ZK3Em5LiN6lY2pRzwI
LMde17zSHNoHJFZ8tyB30K1FJm7aiJykn1A8hfE00+CDrIGwhO+0gPv1hVyFiddEzJqGeykVkEir
hnb4mCALTBB9hytTQkjPdNIU6Qo2t66lQue5HaUSe/10dDNePp9TI8F55foB6mljmwApvgnvk75u
zkgHZaDwvtBBi/pRE8RtjRm/j4uz/XVtiH+azwuBYougwFat6P6lAcN/SmyUh3Q4tbMnemsrLcf3
1/YGIzPSi55Ux5aMeIvwQpmyowNnIoewp5bvxKqUkL/Fysub+evZVWx/QMMqY8RNQ/VQW59IlAN8
NeDrmFNeqM8Y7NZ2M4GcRZh5jbToumsroePnbPRQtDp3cfFx95h/jYRxFJ4iw7A7mv0iGIe2y8Oo
U2qPBA2jfNZv73W/O8aaitJfUkfu2V6y5uqbJKxwlP5Whd+i9yDThvKzp6b5rdNLR1UQIxSIiWCQ
tJXJYVNXsZvJMzX2GWbGtwq+2h7lAT1qPPho4/LKJZ5b6v6llPJaIG1ONSjPwV27AtZtriXX3gUk
QBBs6S7VPOYfEI1L+YfV9y3/nL86jovALQkK3KSklc+Y6h1h39wR+20IgyXgqwUSFX4nCEsv/soI
NjqEb3vEIdfPh9chtd0WeT93gWCfEIsk9y6GHJpBKxlYjONspM7ncV/gOq8q+Nxi3Gf75W9f2XqA
5BeXn9Rj07YOQ1msGrYathLaoDFJ7fJDIAllXLLcJ4AH5SDjKnKGcIZFwOO7rmmVvm3hgrBj2Mh5
L5ySugbisdsWa35g5sssjH00bQBvPHvKDrO9KnNCbjgzj3PxxGnRB+TFViSzauLKLsrX9DX2ZouL
FAiAKVTl4gghxXJoGDgaUZwB3EX7WIdnfhtAf4hivm3yIAZX56WaCEE058ugLBSdvezoLBZra8B3
Ki8xtXfjPi+UwTLZTgCdBDQjhoVv8WOHX8ERAVGe7Hoiv8lJHerujWDyUuUBpU2OlFeDlmGTKb3H
cm+mDjrTvHbVMQkwK1ykUIjKmwNC7GGM0H1taNxZ/N8bSyCBlmNVlMTt611UcExTkiAhHgrLdnoD
pAN88QTK+XXeNsGKLJssJJ5YMG5qkNQtb3HNs7al1hPRHf+966RpBLBHTqfIgCkdbBNKC54lVRMP
2idSrwD5n8/JmF2jg3YuKiawbsF5Qn2WvEt1KrGo0oXKa2R2xrWfZVcuCs5rscgo2NUjhHoqO6kQ
dngVkF0FOgFNLGmHwWR5u1wn65ZGaxE/pX35Hus/LhF84mEFBRhril8GCMxqIHioF4JERAPjP9FZ
QfCB0X8w+U0OaoL1n/2R2/3lMyBWpG2eSbyAxHObet9iczKWk8PXxg2O0hKdalWf3tskhUu5kLFw
hmUhJQrLLdZbTZZpdfYEQ0yl3HgO1K0H5o1fzLGTTvvggrz8VARGGxXOcJtsYf7MXYIrUT4RKKTW
qDsms1eF8PLuN9deVXMZ0i0nMQHLcGBud7unSBVjukJJgKW6guz5nW1iYMXWma5Aam6cFhsU/J6/
0VLgW+Tdyu7ub/wUYzm5M/oXjPvfrKVvolp3eo4idHzaLvyDXphe3BJvdQRujg4FXRrA0g0uzONP
ybJrn9Hab6R/Hpy1gGwYfc1J505gQIPdOBr5jLLS6LYLb8elkSTKHKddDwJ4nQp7QC5Z6JaRpuCT
fCMeI0bMsDN5nSu9Ira+MRGPcpUzi0yGBsJZTe9iMIWfsR+XZbjZq6FWgo3ci/0JdAsIGMs3309y
YpMBUxKFGVlH51Yk7jxET4P5Kq7FkMsSQlbCki/pHCfLuDcpBqufJOWYCopJRB6fkf5uJrrxuZM/
IDDf/HrqyVUntrkALqwDrwIOv5IQwoc/3VvEHKxLz0ZZr4J2Z7daPVvk/Os+18u/nzIX75RTosei
g86cQaC6RXxscQ8AJx/fU1/hg1vliSKnANIpaMwaN6yAe6rrylL8k5xeRan6amg07bkHNikWL+fO
GEb64cw1EmknhapkUD7CmiUFV4f73tNZ5fRcIe1FAvq2wZv7DScW97fFwq+62fMmtL8UpwOg/ZXK
S4+2DtWjAxAqDDPaH0iDJeDayjx+PignhlP0kp3EYSJfG09GEopvH+lYazJ2opkdSWxd7H68ikLF
iCcD3HNIixuTUrXJAP5uXd4Ef7wIg/HBSdyw7aQWq3ciFB7DsiKNH6IUrNNBtF8hkliLIgu6Zt93
h3WS87bE3alx+V7R0zSJEAkcrxxg2AzIqYb+5OIydrc2Np+DcKCN2IDNKATSAAc5wikzV3hu596m
sEzfXEPGP51I5SoYM0rPHN80o0Z9Dxsab6eZBqZTgv1uMbEg26XDg0tgZUC/riDsGMAX9lTUBl0f
72tvKvjsjhqLKqk/6d9EU1s7j2qZeJ55K1LBpp/6KGUIcJTR+u50ysmai5Edhey42FR4ioEf6oqJ
A8l2/7ShDEKDTzngARGcs5nAFQ7+so+cL5jeKAGU1flpofFVufqmySVtcVAfMy1ljBPVBDaNkBAI
K/WcdlFI6D1tf9xpf0MSbZrAgMXWiVN4kenrgqah2tsFcFgMMwI341CilsIdf49f/maIunUWpeuB
rLGj5lojjmqRbl0zMqjC16WXV0FvOja/293ELAyLAuXrkoBAWds4FUC7a6WOdV/GGirlhz3MCRXW
F/7ss8CT81YQANqBExP0sVaw1vv9hXYpyWSWNkyu4qlKQ//gSW07mjypghuhSBYo4Dq3SOLI6YLp
mCgNcWZmBYEUljeB+TaZkGvKSLCQvVCL62VejCpQhki4ltDU/lE4GaS3bEpSIJYT9BT82vVYaaLP
4jLSBEEMae8KGhaDP16H4tlspnjJQyCAOc9d3ZiE86iAiVwtaxGDahGJU/pV8rDkedzMns2HS73F
9vugbVQ3ahmEehIK9QVhWW4ipd2ftJ5jKYGFfimvDZhYQ8OVk4RTJV4DN0tvYYJ0chF7ObaxUGfX
2fBy/3pvABp6eHi9jwwI1LTr9t11UfVUXvJRCB8eK6IO72a+KsuMU23E9W3DY2CH0q5AtGmDYCA7
+yreKvKTrmcz4e7anr92T/N8i/wz2x8cl1C+X9xSy78K0D0KiJLzim/TqS+oDMqR5hGMSF1VfA7L
tkIqvRV8oM9CgqfONsj/0X1Keqe5mRBvFu0EvDnQ4ApDwPMh9keTF+n/d07EZRBX8gfvEatqs/I9
0ikPQEc1cryNsNixExoaCQ2Tq6rI86uT+h5Vfmrl7rFoxI8nfBuAZmQFMXuOazzUf9xGHIeUN3x7
lHr8R0IgJhD+TalWkGLD6hvuKwvlB72+IePKL5ndmBO+LjEZ2fn1CV6VZAnJRuoqmLFayAkG9j3k
iYhVzx26FV1A8nMTV3I4D0xpNIcv9dFQCm/wKxhM6uJejGXLos66k37iJFx97SVL02kDER1caYPE
NdOrbPgpHYG9OAXtP8Hzy/4Tl7Nv811goSz8NdpVrwL652C1rhBj4KxRI3UhE8Htafct6uCSpUQS
jBY9TDPMo20cVHOHOFeMeuHgXKk24FJF7WLBbzkYu/h+w3tZbErNwWS6XJ2lR0Jt0S8m8GTvlZ6R
SF6+NIlDE0G5f3o+CFz/vE2Fsx8rNQo65UW9cHjA2ZAJWIaSHVIE4pDdGRT+07Wjf5+PnRwx7TwW
jWdhcLy+QfnRXoS/JDnagL8upfSEXmXwscCIoKSCcpp+ldk+KENtlD21xFH+7zABDq6VTv6Z4Qlx
yYqYfIHZDMLguVJafUSGujEXvstEbUjDTymX3ks2UBt8TJzNPnMqz8ssEiyCchbnxsIiJNdxJe2L
wT8YCA3K4ibHwADBEu4378GOZHpIeUZqrPsjkg+DS2OE3THScM5XfeVS1CjWeLtOpo+CFw3SSIMH
S04A23CWtCafUY2aVcaj+1d/8YeA1vxBVZN1rMp7TYA6p/mDZiY0+ZvKmZFhmRd6R8DeoJZbNHzB
h1WwyVxl3zDnmyPJ2vfL736qho13tteyO0QWh+xvRJ490SnS3mwQbzvmC16kozXQO/C9KlTa3WjL
m4y/42dq075zjWmWCJTL2dcJbK051b9t9SJ8o4/kEgR20vWHZzOS0NMXvhCz1bXCr3eWLccLxH3I
rqv5hHQCwDZExfH22tmOmadnq9diK+xiVgtTZvBEAHBQVOpam5Qmhoeb0FgJEXYKiR1Er58lqd1x
goeJP4VlOvqR8dvdulW00Q0YLretrYbIZVYZ65EuF73Ol7z3bvHsS1y2EdNpZWjyCCK1SA36+2vX
egwIlx7R9eQi8U1z+gaj9OYDNg11zXB0YX5IWPeUlfmuwoZcCknd9c4d6I3O8aNA37aZ0Ufe3u7r
P0DlS0o2LvN6siNoTqov8kyLZc1X4ifoshGxgzxlEYl1voaEDCc1PQ1++g5SVWJ3JRj6kSVzoID4
qieWgzU6UwAwF42YO5Rpr0AlRUBbI2o0wYZnus/FuxASAQ0BxoqVN96eRYb30ma5RthibHAq0gYN
tzfHXuNw9d3o9Xn/s5dJs80AHvvpVYpA2I0f9ks70TSlCJ1i5HcabSrzn9lgRkbNt6BfvyuVhRi4
g5WAXTDkAUMN/fIwxA6lCeUFH3VOvv/rnhLSH4fcZiwqTl4Ukrpl5iZk8aTywJaWURZtA6pvvbHd
9wauKBjOi2y5VIO1r/zTKIJD7vRRPKtYvzsG2v/hDdvrnS2NUC7DIdDIX/tCehnFPvNLwFr+qN0p
g4bTM+V7oCbj2Jl8iRH/TlG4nYm4Lldk638LBWnMdZfUXmIqenWcRzoyuRogPhbl9T9Ae02IXocS
OGKO+AePSSJUvQEAavlvv5mlvaojYDlFOVFDlo2zlZuPf2LbpW/t7PiDiUnNupTwrgEda6R2gsNh
3g0j9Ve4roIa44g/TspFLGforjoJS2pW7WoTxQ+d/5CWrlTM+IFOwbzWcmTZEiF64ycJ+wNOFuue
dKkQx5E+n6Q/oq10ahmq2Dhanpj1GiRsNAoDptH3Abbp9RCSV2hGLkXDYNfno1UfxH6lwv+zSu7c
bXnrYxdpdpoCR375RnzO5lYyHUx2LuHFuH9mTqwdiY7mOklcN3Sq0q2DavWzgRxMB1AdggAa6MYR
HHkr3EyBVb0nQYs+aM9WhUko/nhgMrlZz2GjiR/vK9kiyta8AHwjWwyvJIK3dPXhqrsVlsz8UeU9
ZgKPJFokVU4mIrbDKka1/HXa8J8YlehuW1gjzBOwIH+VKqbcjYiCyUOjo5NM3c2wvrmYW+knRJR1
Vc6XnsXvzwHcqjgIEr+IeHG/qkxl5d55aORrPBgMvU32taFKhFW+hDDNqeqGn1O/Gxavcv+rXjWI
ZzEPGSsa/BcPdSsWEjriaE6xbfdoWvCvZfdRfb3xjaBJR8OjuBptW2zygMHwjoOAURyR0jhuIOjC
yRh4pSYxrO/0y1nPipEDI4kJ02umaDpv9qRWM6ScTeHFkegOU34LEjvUlIM/epOYvDin+fEj1MVB
X93o0JWcE8rlDND3nDIAFkp1gVesB67MxBmYSVzOgmTYuOlAQ4ixOyjk7Q3ieotuMtZrYz1Iq+Xm
DIhzBpzjGgGSYAfRj/XFE1Xfz35bkIHOmB0wKYfx9poqYRPqkbXL5y5eLlNHQp4mLxUWTynnIbMc
h/TG1FWN2KMru0iB3Vt9FFuigIbZkGbDSWvF65w+/XsI7+ZLONv8FuwmUp6Hi2aYhuSk/piZyVHj
RW7vShAqOeoEi4fduAz//yzCKwCws0ncbspiUQfRWXZWLLgujjgcfVug4OpfUV7fLAkEa45OikPx
yc61S4cZD8mjd5zFH46vDtFLCEZDuD2f53lyAlqxVyqm+w0gNNETvZa3zS1jCwyfd3YTrYxBbjT8
GWFk4B47jgj9gcSOFpqjeS6JNfafyKmURslnBRvDgzUbPlpNOPMV6KvEjGVbkl98z6dST8zsUAdi
W+SALvPkalJThsg5RZNJVNMULVUHhssDFdMYvS86KwK9Y3nhKiHafwWxPPG8qXeWS5gTFot1VudM
5UV9q33niSo9c6YEwVVIdmSOrEPcm7lbrq+bEvmER3ZOnEmG2kOgLONVxSen9Wf4OcVD3ymdDXxy
HkiFbmPaZpjdbZ5pwCY2sFU2rLPO597GqBMQ0sVe+FaSXJBZTjmeJe+VXpuEChhq90Aj8K2mqQn4
X0i+fdEqy9fxJXG918Mo+RQopIc54q3iktZ3eYpOmwO1WL0u78meSgxL8CEVRQPKtEu1UMK/0ROb
qgmrWBB4lPADfXB+HtZENGNnvkqglpknwUiSaZqPCsRaiKwP9i6qYgjjhEtI2KOpbQ2LCL5QHPBu
r0Rf6sBOBWgqJd1pELfeRII3ds4rkkpCWxZ+aZCYxLhO5S/318qhAHN88qxGbW+PgTMCUn6ppq6M
NuxJ58/nsX7tElNKbaiEEnW+9YNBLZtzI6U+xMt9i99NHM3/yMPrm55ytsKE1o5fELfWTB3uL5J0
Rs3NoGxmbjTWwKy7ozY01lEOmUU/aIuVZBp9IEq4AigLUoZdOSlMno/9gRj6h7KIDxeXQ3o7a/EK
y1F66VAcUFB/lGdGYWbPGD/135kMBmVBZaDiyiawlV4xcCkABdGl+zRiEurxAszUxu2dh9ZuLfC/
TkHHQMiVFjlcYQWdzqDTAjGvs/KjYZKC4cAi6k2DewZb6wst+NEmBs4qVT12ZqojhZ7+nvcTItuI
pyMZnEmUf9dfToF0K1bgdU+E6JPA8veNA8N8QNSoqAfa+vxxYo8EtTibdN6bRKot7tVhge49Htdt
ysCNlE5ulixpLmwF1jXuy1o3oqg8YccMCPMaHMLsCb9kzInaeo2bW6idhlR7AqXv2oihlj+E0qdP
Zl9CvMNIwsKUxG8SSaaH/xM31JrUMaNjZlZv3SObGSpuN5bbSC2eMqZUKibv8mndi/KxQxDu6mrj
7yKqUsVId3r63rm0wz/NzdlSRKX8G+7/p+KLsOg86Jxfiu9QMmTUHZ9doqXaETGPvs/ztmJJjufP
0M+91bY8xm1QweVk6kpEJx/Kzdy9qfBhQ+iLuyGeeyyxqLqMPjDDbAroq6nB9RTHRa5QxI3ClGSw
rb+WZC8egI6UKVDmN+koIu+y5g6Zlb7aAk4h3NjJ6/H7m27tjzVLqUhIzN7XmxLe9zTx3GDSbQ5H
ineAaIjNAEayN5AH9ZnIt4sPCd6urpyd/axlCBU4Yn3hufGrwrQWMP5XaKxYCkZ0w/fagnlJoptA
vlL7ln57Cpr1WgeR+CnbUtnEdzRpK1OHoLa8iM3PtVCi324iQRzsyYM5dq52dlCrTmikTEqykjlh
9eMgZQQRQLJOLyUhih6DPW935M+FmN8b43rJ9yfKx9wmZou/q5EUvuZ0ACZc1DEZlTvdIaP3hDWS
OnpKZ9omRaJxaa8jdWpWIaylpsEawEaqgQMXmqpBBJer72rcXFc8HlbE/lHGHTzAtyVMKuMil6um
HzrplFb0R5aKuepsUSzxg1UxaZ2I2RgYHfFiCuQwQzwUrgeEhhkMUrpQEmAeYuQAoC2U6DiCMa/A
vNLjSFxnUNvuFizTh3Kfah//RRrZCjnggnAFDI2e7XURCtDW+xJFWZp8Vp7AYkheMwE/uOooel2t
HCTS57qfyXLCmKcZg7mpk3g72FRNOyM8yR6Ux/Kbayw1xBVdBSJcQUm0JRVZ6Rph442krlaib05e
4TCtpoLO+o8pPVyxRK2sC9yhPuSMyNJkAKgFG2/qP+NKQpQBsghwPibqZbHB6Ngh/pU/YHHlUgqa
qffVVGpnAE7YyfAmfFLfAeWN8fBUzP6JxQUjUEBoJHOXKCrXbmWroMTjuP7uC712y7WSEwi8EZeC
FryzUmni6kJeaItxxo0x1L4tCXIFcXbaAycogtRE6kLoVOGqAForUO58Z89aGx6XOe2jHo63ppp5
BLdINgOZYuMK8phstK5SfGjYxyG9250aVkRk1tI35JImFtLf5SkhsYMS+J2K72PrhTu6nUjhz/U4
QOrW+MB8i+6G+ZAF7NHmX1l1Nb8MnRG10OJUK0BWqjejFtIomwwnvFrw79vn/v2pu/NzpHWitxoA
OfXFGp2SY4E/4phpuv3PZNu1S2BKtNRNGMH4126wOhbTtjULAk9kxbVMiZxtqsFjs3rcYDu1Ky9S
fxRfplvlFr0U9PaVIt8dIM5OHB3HpE3VtY7f4vefFVufiD5Ft89T28qXGnvh200L78ewMChk2pR1
BINfipivVRhpsRNO16Ot61b/c0TA/QQablFAlz6mZwPrsYO5o1hNHSy629piiIuF45ZG17RBYovC
vFLBJNW06pEi0EL+H1sXaMEIHQz0ROl6gcJC1w1bTGVvamSqMZPIKpzrU/vgKPKyyEE7grTPuuML
wl8hLD/Hl2dPuiKYk1gpCyU84P7xmWPfkEnixjeTxo/BzEZodIaCsWuegXHpbhMOx/+qPjuTSeCY
+wICNG4H/LjSHbykefmE7OxqXQevBtyOc6zBG9rQDB7+XzVpPHzsHm0KM8jhCCbjy4y+u/61Yndh
ejcgtoQq9iLjXc9pm+2pDgIykjsCRmCD54ptJjTgcTmgDOqd6Tj9U3voACrOj0QryjydW3LQN6eI
leBngRiZeAmHFXT3roXVx7oCKbrbbdkGoVnNzheJ4bPlRdcMOL67e/J4u4YAf8upvg//qzVEj7Lt
qt7tHT1472zAsfvXPPxKkDHbuprjaaAMhMeSxa/3tQtmtYkmb6vMdkYbVL/0owPDCcixhdTPCS0S
F5avAsjiwKSD3XnncevOm49k81w7LUnIbNp2wo0rBzvNhOHY2TDdceVWzf0FQeC8BI5YHH2Ir7HH
cV8wYNw+thf7Wf27Y/29T1wbnL80LCtzgujWOMMI2asDuMU5O72u0nkFkJerYdavQvOzwcMz95Hs
JNtnsGYVrnzsdYE7kaXXbqbJjaeHAbmJTpi6KnU9snYuY26S0ofq3dxWUPLhTwow5G0qKwhSMjlx
+/AXSIkZZCulMhkDgcKwuCAcVUMuXTgBf6ZhenKFVlZydTeH64zLLgqtCInwboFBcDjcdMQaFY6O
onlydeLfnONNXNohkrU2i4IOkkOBQ0j4z/qz3fTnY6xLlOXUWfnXu/+WuDRxpv99dU8F4fhV1cr8
SRw55MWBYjFAQ8xNtShmvztb+1pF+d1GsaMtc2X7+0COS+ZMhPoXLw7LZ+3QVjm91tmEhW0DL0Zp
xVoVu0y1vPhBQEAyoULzJn235IvoXOWNR2itYAE4woefa0Mf3MHZr7FvkxoSVzTRQ5g6+r9v86wY
fsl2mX1HSvCtbcSOToLTwmwRUUjGVqD2KACyrkinFmDSp/+blTXNT/CE4G5q3QjVsPF7gSYEaqhm
sQIwTYBDwKw8xs7anxC3gGzmFwmcWTRyfaaik9BmuhYhdVQOk8hS78GfTSvIgUYNKjSLRmb33Mfi
jz60md5kEMKhI4y6y9XtNmIlAOzgCgMd1gPKoIagzb3AXHnBWy6tfzJ8kslvtjTdV3GaQpnOYgac
e2Ve7UptL+U7cpA2Ftmxxiap9v5EAr1EXVAvEp9e6nuPMGeovMuJPVGn/S8zpNCxGpbHd+G5xmQl
3+7DGwsgqIPw6h7BrN8AhgadeEEwTeivLjr8XdkWTHnQ3pgy3p2Iojb1N6EVw2EBFNB7lvNi8qZx
aL6AQnaLfKrDo5Pf15RHNs4GJkbr+/k51qrP1s7YyAyQUd9m50wBF0vwTrtsi/OG5ft/bspXHu/K
rDZQP72dTbhRbMzUz8W9lJnAIQM+/0gSaoBjo/dW9M8qmT0UhV5aKOkEP8aJrP84K1LmjntgYSa6
5cPi1EQj0Oe85oOgEgHAsggoc2gKnGLT1QXakOq8LJyFAqqO8iYTGlAiXxFFr51IltSzzpF6gzM2
e3+a1p9yd51u4+51qEUHUXdz9x/66E/sKHSoA2D09fAMHtKAWGKLkytHUNMAT7ORPEZAqc6EXehq
VQGdRMxIlAv3Th0wt5W26mfLLTGpGXgGhOpQXPwl/BKPF779lFa6P5Cm0kda3iZZuiqh6N7jm3fq
fxwhmsrIVTZm3X5WXYERWBQd7wtVsgKQwipkOSVqMCs1bJR4+DVT/NCl/De3rJDiT+MSk8klPvnf
dFiKfPpRfLCUb52hTreQPWaswz2RIh35smIQkwp+rGukEOfujwFqysItcTl8I582hhkvp3AilX8V
+WpalLPU209pyr6aLg56TVop1eRSNN5KgAfCJ2ul+u1fx+9uOw/IxzqGBHvj19IDUg3/uF88n3Es
8dsIn1P954mgoyuJ7Fv4CG55+wO14LdiIum1sd4Ca2pgsi94EIMoOBo+l+vQhSbrb6CuaVQyC114
uLNZrc36gAWM3i1LHEyT+YGkKtZM4yTvkzpngoPJixq78sf/4DrbHbrZwmFna6O47biG+ipUMevl
3Xhwn9eik9N3YNzq0GpX0H8PYenRZPs6nLq5uzfx3aipBSLoZ37xypO+wytG0sPpJ26Xug5ur7E8
N+8Kz2jPtd/muaO3zBNQ7abwinshRg8pIdr6ALNptMmzKHijiho7vZ+HrJZLYPHUrlG9wp5+/FEm
/YL9qdeQgyGyj5YYSQbM9RwiDcNiFTmvWovx1ZuykYpaySZH+ZHkrJamQiZwXo4l5SeMgRcCZjdK
o4uGmVbk2v1O7MFGhDktN6uyG3T64BDdUF/pSkCUW8oEfYuYyI8SfT/EZh7MMRDEsMu/6eKMkl8T
5YG7PPrKO+rF7xgWv636jw5m4HXkEmT5Ftq8KuxrPyrOPsjFA/Tclqa+U3XBSE0vAjOgVDIQ6a6T
lCpT+iDaGAnzwKS7BYR+g23LKh+JdCyM/H4e9HAQKL+5pfpryR9E5u8k6dbhpgy4GBNpDuji+8oz
jaSx8N1pLD2eM+LW7jTDB06rQnwwHreel6maf49vws+QSTvtRJp1r4wzUy/4dXR/BSKVfGcVE2k8
aa7v840/XoGL++JHVxa4UhtSZ4m6fO8mUiLai3QhXmVMhcjCVWAZyj4mWrwnfSuV7+TCjCGaszBf
D/1dqR02jzm1cD4YMilz8LE7j5NIDDIF2Fqqhaeenz8dzNRp9+Au9MzFFYVBg6YoXkjqNiXJ9o2m
Mp7QOnfzPgi4ZhwbRuBGxVn6qeL1YIyr4cIesU7JXsaz/LjB+EM+Tu4wz6Ak4m9PDE3EIi2UzMHX
35WyrSStpYEtW9WO7YOVy3ZcBfSWpLrhuPiQ1EKRU5KnCZWoq/1zN/i297Wr6jvsduBXJax9xriA
wDe1RMZ9vid1a5c95uBNZ6G96Izq5QJCGR30aK+ZnrbcfzCjLWlkOb6VqXht6cRZyHVG7b1QCsaI
QDxgfmE1P5ByFbr9+kt8aPTeAKhsuX2OU4gHyY27NltZEO/n1MDZyky0Q4cUEVxpDb6OSll5+/Xq
a+pM2Jr2I/Xm/LZdusAtbpx9jLSz2L1cJj9NioIGAkLQ2fdchfqEFAfMde3zk7GT0daaZiMN32xg
xUwW5HOoc1/cwZ70z3g5K3r2vl8XYGvjAzC8ahcxfsPMyHHp62AgJYnphMGK0seNS2i4HW1hIdUV
n3THjiErU3mxotsme1GuokehW1HpQsbwFg5HVZzo/XB4OYdnYkKumHx2dYsF+3VVg8eDKo0Q+2KY
hlSYuBbiUzwX16e2driHyxzDXkqge08XYI1qLLeb1CYmR7YTLgsH5Duf5rzXUUIxpBira8u/3d3m
Bl3rxScsuTO5mC7TwClzsELGhSAICCL2qUWzLVobFr4yagyky20BdDcce4AbLbdlkWQZQc8dJeqV
D+PjVauGvo7VybzK1tnhZ2iwl42k19GgamQw+ohN5xv0IItb/UNIbi6V1LHzSJ+MPgXbDOZsVxAL
7wGNvDQtgT4sqDkA6nfwfBUFcPjyTcdqUUHExxOUZ0z7eD3qIFBka526m06XF7DV4Kj3Jld6nFom
A4OPdPYBjuUOCZ3gDHB8ds4W3GM6UbQd1sYdwuXsZjkc3YKqWEocvlJbIjeIzQEnzU+9nEifLJZT
7Z8hKgUNQ1bQO3e4jIAdSeJ0SB/EA1vbFfXbN1mDjKZ5RsgYlFyotKcapaTtXlxzkXs/Za2JWkGp
y8JWZl+kqY7hSMfhMr1yp+VPTCfgrXJF5EWQIdFk4dIiCDoFdDP6xairUx8sf+bMz8qUbSkzQbD6
uED8EQMgEPB+giZQkBEMQGgD7sWABTq51DCP7jsE+benBYUmCGP9s4tYeSHqQdrySELdUo1lzyO3
OZzVGbfbIVczO7subsnwIGYZSRhSoF8zSJHQer3umd9ovuR+bwGSbgmcAu+yfNlAVf4IpvDXiDPs
r2Up8NCf3KKCoVLQUWXrxNDQsXfHxvriIvypqjec3DgLMa1q/pRFNYmA+kY+FMuUEFazqfPmA/93
tyHI8PrZcnTnPIsif5ot90bMjlfyk89BAHnxbKiy385iy++FQUNvBz7iNa+dLlyYORE0eWzO43sW
BzF8dGa1ZQHLRxha+n4S9B/5qpz3KL/ANhJObfHsTYOpuFDwBLYMltNWOaCoMXAMOPBIa1fjsbzN
+rxhxorGCjfv7tUOaKaOAboxpkMiIyo63EXOHesK2QD4SCz9Kb/YOBVg/3GaoG9hqIoSJ+Ii6dRP
rqgKycp4RCoRf7mhuf18gPymOk7DgMwbJMVzAynQ3ku+L0Bo1Y7J729i/58+xZO4Hly3Hoz8IaZ4
Bv+MOnZ+70V2ah9Jw1Im00oCrgTRpDYs2lCcfjNVUcNpZyHXTaI52kS0S/sunx/xRMTEexeUgGFX
jpQFTPZerZBGmQDTNOvtfD0VuxnAnqlQ8OSz5jz15eaGgzpufrcTTI8AV/+1UC0tN/Okku2wYtRp
brfEZHToICEZ1ssoZlaypOGCvxeqDrF0dB1/FHsX70YGfneNOLZXeEeIAKDcvDxSVj6Ii9+fLaGQ
mfH48AbzKHKLCFdcFDQvW1BFEvDpOlZuctWlBRekSXptl6zFgV+0SNk8vNeqoU4k/IwoQ+7Uy3gi
wdkdSWGAIUKGPoQVMykf4aeYbxgyIqDD5YuvRgvRgnHcjJwhCQqY4o30OfEqC3szFkPfShKCsyCP
SBXGj7vZTulzl6yZuyle8w9jtNNPpNFCrJ3/zsEE1GUA+1vDTBs1hKPmpUqEd3Kmx2DvY/9FGNFH
BX/CApigqYgQvToplnykBeqX9D+2gV2LbQJorWbFvtqf+zCLZNph62+OaAG8kC13UT7GUZhVWiPn
QZ54Mo4fTq7LFC5OrW5zYkT99My9APaVggtX3rWTtr2ezHspXr+Sda9zZ5O8SjV3BxUrgNM711x0
5vXNNRKcGLgXDrs46s5KgESkSl5DY+W0aKOQVsrJ9c8CjtHoMI+tUt9BJXC6l7L7fcaLpF3S4WhF
GPBMMZCx22+ugCJVF/1w5tPNHcelhx1x15mygoquRjMAA64RoTN3nleEahPRr9IbFf3obyodtzKB
ZcTix3NVP0Wae0maoBV5amFukXJN42W/hw3ZQfZM/lQyL+zrLucD72fx9yA9xrHDSS45TTDVFAEO
a9cI2WPRpj/toJ9qO1kU+wmC3UPiJ1NW9Ym61d1YQcNbb8R7J3XHdZeRM6DJzuuPpJa5eSBrkt9g
EWTCizhQp7pvZZNTexHwl+0QQa/XTOW/MuPD9OCk2BWcrJPxclwECDeunkFmwkc9l/wtzd1DlHwz
WCzPOWCOlvE2/ELYCMEhpabiv6/QTtpuhF4MYBfkkJfYuwoJ/my8L00uakY5eySYgb6GR9bPNhu/
LpbVDkPtICawNFcwcJrz6gR02Zin91AR34yjpxm0CCR3XXFGz1qkjKHvdHerLZ6vTonPDMfNPbm9
zZnqHIJuyZd8mc4FoGrlKrTy5fApVsnKSeZcLAWdi7GRlAifHjJ4jccbI9ltKC+obf0FVZ43MyO5
CQ4VKTNOkx0A9811NiIRNsgAIX7Nv6Cfr4QI3iHmWZoBYG7/yjpvfI2f2L4K82x4d2Kewa7iB11B
LodCvIfC+zqBEosFw0exC4BCoBcAby7Qcf2b5WRmj1WrPVUOfNRMG8Iq3XOh+zI4byBs2hWbdVTn
3WkBQrlkjI4kfkWxI5rk0vq+vHT04rghVtdR6E7GnnaNpfmCR/vK0bHyLzfea4xruodwqtSMYae+
+sa+PP+JAVAzGRw1ynXmk0JvNlgitf0lIbzqq6coVmzVh0Kw3qMcY5abyD1MVyF7IMQhqRZSanll
f+yAKQECZ+JotbSWrrCa9mLGxVsM0m3VKXtI64r45ws7eYJOUnsC9KKPw/F9IvpffZEwGlLafxMj
rwSJ7EpvjBrrct7Alcth5ldH2iLOcfribpbqg5SDEBOrrM68WOU05Yca+GQMH7J86vzdTTRPk1Ep
ACrg++JPX/F+nKJYgnGlBKUD6WFzdHDFeByRcG5YWdn3M5LbDAxr/utgOaQ68yEnFdX8yYiHGJDX
PI1BqoQ2Cvwrk6LqC8CDVxBy4IKh6eBPdffcAjOb7ZoTw5nwvK6bcQNuQZq6tfUsXuAQtZOsi/Gd
TgTeaee1/sIIMKmAeptRZL5JxO5VbWi2yyftdVPjCawFX933yuYskAk+69USpzvrVG/3B0lejvkN
akeyghqwMOeNQsQDcojJOamz+J0NZ9H92rD/BWm4fArvDde2Z85X0QK76+/WZYtSWKZpT6/tKJ6s
rUrLAYaYIsQe+CEN+8A+UYdoG+lLotpFAGxcKOxvCznSB1A5hTEWKhaDNh+Kld75MtvDnZsoe+Ab
VS2Jf1bnaGVO4XCWPQDtS2afornXuPdBj87YVE6bspRfCNT+Z35ZHdjRdyWNjbD2WssVN3bZcSYT
MWGUO6ijpKGcIWcdJVZKQawH/dd09u+Ed0ptIxwjLoJblcrhyVzUOKbZfS/N+d4Iz3aXvnvcZROL
wqg7flrM5WlgLBEJTzUaXsCYAPCU0ZCDwc6tmr94XUFGk6fUOzc4PQMXMNtzp5m3zgbYDKpBLU7x
Z6dRXKXCAijA8SiaGvA+CiueFao1+VamlHsY/Jl2H33RSU5ZrHyUU7lIvDe5dlYNQKcvZhtBcz9F
QyD5oaXnLaCzMraAMJBFF5Db8AMxYYZElC8smFH61hjdKCvpslaWb5B59DqgaA4tIE9tKhSbbyze
N6uj/95KfHZYVa+FYfVvS4bqfQj3QUNcSpKFTNeSrurshR7BzUGOsmmQTrpopvMwmd2twUHh92c9
65WL8XYrH+Fjd1qVyIEen6FJDPH3B74VehRL2oLOiek6avfvTr4qJ8J75SdGpJwuQ/8m3Rr8TXCS
I8QlY4jfxBbzU+a3QwqJ+3h2rbE8/9Tt0ftLPfRKxaq1HR3/iq24hVYqRsK+Ep4BIeSiBpT7ZhVC
xddY9VK51lyRnFGIXgv96KqIocxFUGJxOlvx504fgp3VvdEAvwD5jSvmsXFUvOzkKRSL2rwaoaao
r1zKi0TTyJ3crBRkwCREILCzgmgsp9rVh+6UdgSbYEklOvoJw06OQrWf4JPLyWAFawxIFo/SxxpC
E+hMtlR3Tkv9Nd3IAl/hpeiHchwAw06h+cXkjggW0vsG0t2dG5uBVb+9y4xXtafmDd4ZlEx01Zyq
mDBnvKzR/PtYSUzBpaW8p4ehA5IXE51hD79ccDO6J3dtvtLYlZDVOu9/IqibxsNEaCzWgrpGLiWq
D6JkilDBC0MMt4DmlAdWqMg/duyyWZ4Rpqq9azrmeMZ+UGagJdP7ZJecYTbaHWjB7RS0zq+Gy9Ew
23xHENJQsPao4wC1nEU+vOJnuxFXMgrsCQdKbTF9OOY9MCx1eIfiSVHjXNA30jtDLB4mpptlTx9d
NnWWgpLIPZG3PfhDGfooA9VGBUyIOPl/aR51mkCjSVNyWu68q64m2tgD6KynSu7nUs5VopqN7bVR
+4yTs0WIMAaD1gNAxPzUshZVRDDn2i9af9T6oDShDYbXUbN1MUtRlRC/OWwbxa4PsqGqJ+IYcLMw
1XYgij3DasKJNjbbNh5v6RFe1iovQ9hr7Y7UdZijieo93rV9KLMSSgm8BFyAtoA/sB0+B0LpARQ/
PYM68rvsZNCfflv/sfCT1RT9zVvTL1R6jjFlds9vMe2IOpqWwzpyoS1PAT/HOvFMZBZlbkJs+tcm
N/pdUFdF264WAMP2Voy1kG6qjR6MqW5XkePflI/lP6qr6FWu4QytoqJ/uYr3czOJaCP6f2wtQfpN
DniyD2MHZvI8rG7Zq3J/FqqLIE7Gz0Tb5sQaV0bTfHnNJ/AJ1SpE5LaN9oHzMFFau6SOqG1xf+83
XFILAfjUEXKehtR5u5FxbaS6PnQi5Gb2ZuCMQJ0gizUnpXQJtfcL42iVBmJbf/Us8QzeV7AbCTxB
d4RhRmOsE6F0P5BM/wtX31Hev+Tr1by1Z4MUc+XpOZyjJW/ifA5x041s3Mf3O8OY0cMUA3CxaoK7
yFn4vUc2A9cOEnO0oToPP0vAvYxgZUqnX8MjMTwgMLOprBe1GrZ7IL0FEzyLDiI2bffp5K7dEsvc
Lbxx1fmZH75mfUPJUaN7HL0IjOhpq5Y2wU6Gc8HmWbRLXlGVmRMekFmxXkdvHo+gnzUd70Pni0oX
Aj/FO6s0la66XJE4RbmmZwdAJSILOi8rP3If+DZHq43Ymrvt/QNL02e/7uBEEJVSDsCkU80T9NMm
PmLCpO1JxBTrxcZz12EXA+yhEkTGOSmn4E/O7qF1MnJWXE5FE2p1l8F57aNESKuI7FJpqKX5jXs6
iKwPObjBX0esKwu+LUrLPuHxMeq3U3Rm446z01GcPVhDhoqDkhPy9TGUBfsUMnj3qkMpZACH9/RK
E3YOPll5ZCaGlXW822fwBtbajai+4YaLWSv7m5weC1waEdjcszA3VrspfXo2/kIEaK0sBw1v2j3d
w82NJWvRq3wSt8FmrSpOOhTO8MVWJHAoRG4LAwFrOCjDMKVFI3B3aKbQkOH6aHufQVdq1+lN/1S6
DOd/0n1ZxtfJGQwW2c1Ca+ieI/CWfOxr4G9xqvKlFPPp9yNNP4ogxMLJTUYbrH5G7TzVFquzYXwd
APM6myQs4cKwyXm5nol2EhFagwtpIiz+to0ytqVgFHfABB/zi1Ovu1q4ixuKadITs7Wx1TDst9oL
pziAzYpMxwPf/Ux9vEkPEx/AcyXdxagg/Dygix+M6SM5gyi3XXZOUJDhMGdKn+D8qg7djuDFU8n6
/9rFZLbIyrt9V9vfkC1U8Cp9ceCWz0/EYCIyR+kTEAmZK/zjtuT0FNvb9fpAtAvQJGY4sVSuqLR6
da5ov/EKNh1Kz+/Tu9AJbazBcWyZ2uo8PeKlbZDn8udI1Jz+ZxLEeoH3brETu8wN6aSiCUBihahb
r7ApDu56MSoJ3sZzLbEWVrnxW04Fnnx+CYu9Ee1GFL6CSStGSk5hU9xhCxf89tfdXcH8OoSFvFyT
QxiKI+mBaXRhgj5EnKVk8LkhiIPQA8GGPRb9JCTGqciGE368bKGCzx0sLky2YZ/QqTFGL9rsx7hy
FEFl4CQY2meYfqKCr81xQpE/mrTzZL2zxf+a3suDo1I6+jLktswf2eikmvleXK1OOjYoJagVTmOJ
h2jSIdTb3Zcg+xytrtGzd4gYe+lvupaB0vApKuCzLiaTKdElSqWEBAwJ9hW8Ta/gMXMUXPMBbDXt
1sKOBZrEA5M9yZklSMMeC9gpfa7Dr7OV99FIQQUdDiHW37hfWQ5U6hHan9bZMNWDhu2AFTxmDAFh
ZsxdNDxyc/IR1GHoVwalbonNYfr8q/qNH2XWLBJi90DDwGHpl2Z1mRnrpWkBebg2vNF/NoQYIX7K
wOhgkvD0CRh/dXpfXc/TXxdI3YJvdxEcizeqYMCTdmptNolQ5gaGhrvyG0zNMeaDf5U/6LoiHM91
Kq12J3AQ15SYEzV9Dc9UG/uhqlzjDVY2cLn0evn/yZwEc+DeP43XmI9sjpcpgGj3hz5uoMnYJPX8
3NCh1KPSlfFY9EhwSSJIhJPwIzEVTLTuu92wQcmG3fE5Oxf3z8M73svbs3uVEo8cnHO3FdVcbUn6
VaFsiccBD853Y/GHbqaczuFq/kGlrJwfu9jQwV9ztaVxAz+h1W1TEeGTupjRxyfYoHBGpj2xR7Dr
woKot6VuEE3tBwsJljIyVlv0/lQBZrxK7qIbnQG4wi1h1S4E0VXVNjojfUDgRF+B6o2Igqtg5RX/
hI2fx5t4pMFV2cUeVUOJdwt9F2b5jDci92LUrEdu5LKKYEwOEKyPTiu95hUQSUQZMogE5DKUhwUu
3Jw0FHjs+NMSZ8qz15WsZhMu1NYBKaeFaxuFxXYC7e4yN/vQmtikeKrhYhVkbC1n0FclcwzZ29zH
aGlHsF87ejLx1kLooXccJ2XcKFgvtEFqRi8ORBQ15udkIMnXayIeNRqpMLGZxIJlYUMzfsr6Z91b
SRc3mzF2pcfn95BGykI4+BdEPs3ZHZFNFRJtXvH25g9jPHLgTASVBLK6rfPxSYzXiHmceQ8qPUQ1
wsROQjGOup4d1leND2lMLEcVqcR8GCmSsD+nzSsQRl02TNdK3MxB1vKQJ37NT8b1lE7yGW37dEcP
3krnQ3M3/6nfA3jgzcpUv7y2DrVAztO5aOxUC7oqLqy9I+lTeApfVonXzj+QeAACTf+vcE5Mqnr4
fYbe7LKCJPVTWACgt5MO4s+qT5Xo9QUyKSBmJBwiYI02lz7yc143iofNXr47Py8rkXc/N/rPcrxv
DzwtKCht7NEF/r5nEZR5v1MkmDa62qksVR+oJzLtuC1026C4TaQhj2V9e+/uZacBKxlHPRN/UNBS
zJMJJZf5SpeN52+DY4PK7A2CehnODOerYSiAjWzGkQRTZExyKqdRMJsryrmjRHwgJoIDP+tKiibR
+QElOdAddQspj5GABtXqGPl1hZayYdCq7QmElP9ngL4ftZTUFPjwbFK3cBpb+OB22hNNzVOmK/tG
/U2uzsgZpSLW1Z4t59thRjtHHKry7p/1z/5itsVoDbp9uYrzsibSn5UF8dmfhOaw8qXnhtklhoFf
dDF40wgIn4msawQe5xzksS3aeyqgOVQqTtai094q8r4NL0mYTqczWkT1prKyu6mcTmzzZiestAW6
xm757XWYL2faqoAv5as1ZL3HH9Z3SvZANiVx/W/QDuNHwhF07gxHBGBPO40HbExRJZjmpP2VKtfS
CdBDVtsVFVijOxAE2wd645r8Y6yNoCoaAYsJDrHoSsDTHfPfw+pRKkIlv3FTKbsZg6WE57FLt2Sq
1hbVy5VGjfG+0Kqwt/2oRTmgSLYyVuQmtzjiMqouvr9kv7+uPEFWEsWQPetWtXPBTW6njLT7MDDw
kvjo42gSODepJdmPSLBiDDjgu+DxUE6LWLiqt63mHdBGNQ3t+Obj8fHKfBQHHieGQbso0KubhBT/
kzpbhsG/RwvYQ9mxondUE/MGwga9gc1Nz1sOQEnBlhFb+CFqoOva2jFO2MsmMGUuwwpVQwQewgqQ
vsvpT1Al65bCIIaN4gy4ogUk6E83Panb0EYYpPUH+4k/ljA83mfGuC9xByZj38bCUgt9oE16BkIo
MLu2PDiZv/3bPb2LBoVDSe0csedkf1BFaKIB6UpXWnk/AXdi4FumZR5lYun6PQeWiXc0OswNl/P5
faYGAPS9q5nZiD1uL6/qklnpMh9Nor7XSGYOT8hbL/gXGKJLvph71zBGettn4Sh6ebyTeg04uMbe
6WjabKw5zRfswHZ9q/1b9MPbHkqaMFGeiTSgngMgMM9dLavCjeRxQ/bHIHMyMKm1ElAz6Heh6kIW
cgGPTt8Uh66QkuqFyr/PR+ThjcI9yr/cJH8+1TYwIP/I1jAUaWSbE/TxbdsCuXynpg3xFD1csCot
3OUhlWqFB8Z4ITMoOW05f9urs/i72EhfOCWqI24OehEbft2/EDMv6nlaXY64CGKi27oI4ARlD/CU
RCoKWcOGfLyXMnsan1pdSpGdm313sbe176ESDZ+Ag7tMD9QLwYpKLXfrA9EbVjs0S3NzVjhx2+SF
GYfGkNfQXXeQRieB2ap2U6+RmhL0dB3S8fL6LnAdQGZkNhFGmfvh4PBNISIUh/kGzv5vdEckq7e3
Gzq2B5DwejZYZuAljhmut3IHTkfp/TWbt1NrdpMnN+mnPOL2Z/6a+VfERuyVffvGABOUF5qTY5Lp
pbGZ8D5Wt9XknJUv+x2x/hXhmGNw8mS6Qw8UguCDEJBnuDubqK05h6PS7F22l1lmAh9NixOZpqze
s4yVugex+D9dIHy0g0hx2UQyKCihvdbOQORRCrGu7ls1vBZ14il22UINfYimuQ3kg3JJOcHn6bZt
49pb+ix5SBiPx8eAHySH/+Ct/d88yDhVU/m4aiaY3Q4L0EwbNCn/Njnsf2ycxQDOsv80b8dYZJWy
sMHSXtLPpRJrgeHKam3k3twWQpbeaK8T7JBsWkk8Wyi0wyMgOLlKvF3qzRffrwxZz/jQFDgK5CDs
PTdC/Nvag0DaQ+utfLHVc63yftYqLIKbPDtVAMIjWl6uxXoVWlXlq/X8HfjIwlxxCVGM4LaAHCqZ
Xjoo7Po011cCsOp4HINBFsynZMnCq1ctLAQ/L1mcqo5GjmWZeNiml3WdEA4jT9E7g7YDfZnGtiRM
tjo97/BTeONH0GVwJygDxvwGFqpjTI/klCoV6SBCAXdNjnlqw6OVKgb24h4DOyff6wmWt5YeHgvQ
rPs/pR8QpKpwKq0CPnT2SeUk/Xa8/LHaPwU/ICtmK3Qe8a/EGZSV15W+xypNrP6Dirn214jeStpD
MPQVcpVSAjSNaafavvhmziWnMmaW5Lc1But+7wTHus2rjb7/6/BN5POqWuNdnzXh1AtnKoZ56akZ
7UeXTXX1d0xNBxEQItsZeTbs0Y9ht87T4Di4jKiXFC1aTmeQBQnlEJgPr36itkA7CUCOoUAxytie
esuSEGtzNmW51qv/V7p278lkx5kB5ImYOW0YIKOQ9+GFC8t9Ee/rLNJrSkoAKvfiKPacyfMJuqih
p9v+3+F1exGpequnuragJmQenTJBqIHE2NzNVXKCavUZJqcUntxhos0WG2DeajGU/t+RjM1DKJBV
c0nCLAS+94lV5T8nBKbYG1BKClYGTmvS+jOzDyZDXUKWRkJFuKp2HPBFug8QHjSGQ6VNy/dJMnJ1
5Y6MvRZ8CMK3g9Tay6BzhsoS4Lknj7/s/3ao2cicBCAdw+xXIhCnAYhilW1h+LQA7zNJxcD/mHVX
MRxBZrZol9M9c9SvXE8govAnK76Uh72jYetbIUOTP8bLlhnMUD1/SfyR/Cvn9EvLGDWagroMtdpy
u08/wW5vFngvxO7hbaCUrB/pq4Uy/eq9xOuAHsitT+qQiAwB4x5XvUp6VRgirLOaXom3tn29tLsC
xKUKNwZPByzjiZtnqq+Q/qd9RTNORUH/7gL12SDXlXLMOSioqN61ym2mDfre5/1pltVwNsh7Tc0y
iNhHFqDg1eTVATOpstt6wK55Vmd5Lr/wvP43rpNjYIoZFTfUNNAx/8K8Q/bMQ80vumCcUMo0beaq
HqUZAqnaswTpcBARaN32gH02JbwnkBy1MTa8FPnY0k9SV29lMksD1ZtMEz1nU3VZ7ygV2EG2ChKe
3FdDXMER2V49HUcNFv5nRrKi35odN0eCkmJkwrGua9T3MGMk80ZY8CS8eaMTU1m6qY4ihVB3jGQI
58syP5hIbuh+sbdHyDQmTYRwJVTgr40u3+6wToI+Wvy+5abBfBgPPE1yxfCOzdrXnWEgKzjBbLyN
RfqcTsNCCXGbv7cRnEiH8BmW8XBSgSyogPvTGiEWz/r0ytXhyTP/4U1J024jti2S4l/gT3jn5wGf
AByMu2LbflWLkjpw3WZ+HapCrUIxS5qwrf6EjmZNHOiF5u/f/3MWZHncEg4MzLSQd5+TtA2H50cq
s4GEX5KL6Y2dMZDYX05ni1f9rPIo73F4lMj0dqErt7oci6p2ltpz2UxypR9t1TmhAySbS0902bNy
s0exN+/KRXpK9wV7bb2XvaPYWvFzJBzkBBnHuq6SuRso3ePgB5+F9gNoNYPE46Zbbi5jrWc5ARfQ
hK4NZWSUv5OWJoXEwHR/O18Ky9MDAyt+xubcOy+8WnpquemfMoVbOhKASIrxpfsdR5gHAHj/jnKg
yliDGcR57PhmyvyTbTmKs3VM5sHevflXjipjsMG7gRn2aWhC1UvvQJcPcJlUPrAtpoAlluvq7Jyo
XTowT9j5yFbsPtNcpid5EqbUUaCq/8iXyNZ1PV3DBIDBn4zXs7DcUooAIIUA8UeStda6+BSR3Wdt
IWXk/gNT5HTLv9fWPo5pcbhi/0tN2uei233GIPbFrFyEdUW69EXH7Hk4QYpne2g/ruoe4JtkFIht
jeU72BHcxtmijKnruAbzb2RyS0tq/UWu75Y240+uolqXguwD1uiKvOxib9W9p8l82THN+zAfpO1n
Hk3EANf9TxewB+dCyaFnu9kqcmOKUuHYWOxKOFHjUH0RPFj/5dzIDTXHGW6v5E0t0hXjPaICeylK
j9fGEncxz0QKBws3m689XaorvwkVebfp5aq/HVGO1vvTogVAodSk/0UHSeQmj3fpq9Ma3VJhJ5BI
BRJJhXydOj76lotnCeudzBwpibiuP9P8YHtBodEDQL/bNlsrxo2It7zBMnPF1AONmBqUq9nDQrfO
lzZ+PsUW0Ap48yxqUs7PRwkfqDh+wG76/RWCx3R2yhZ/uLcxU3PllMKb5vZPqe0oP7vEIdaKDCov
q88/LaXCB6oic+UE3rINlQ/zHTG3CATn1sxKmC+zxkGfBS20v8AQ1ZM+D4TV/ff9LGJIoe93coCx
maRKos385eo6bCQSaniWa9jzb7rXAGQf6r5/xICHhteLCajQTJbs8qffThtlZJTZ5WTZDNbdE1Ep
braktxClYof7yEQWln/RzOybxQM3GkTvI8SZjcjvE2SbTEN4s3CHTatzuI4eyk1mGZYLdmtG+NG/
rRAM0LCxvEu20HUpJkfAOt33E6gGhD66pid9yjCRa/nX3ymOhkU7SL6iPj+z9qepfDC19KT5HtwS
lFmnEVR49FtRhDXMQ9Okf6m5xOB0V9lOjsEtlEkqLZ6rqCeo61Vk2adM0RtoCHPTRdOvH2q83k7c
LZBsqToE8gnmXx73KXXoe34qYqA1D5XMvktjLz6slwgQliyvKz6diAA99Qrr/MORgc7S3ULkkI4t
VESgAMEOq8GMMS98PyPST2wjHtvMVJoCpGL/Gh5krBWp4m1F/nLlJH3RD5kFWUbLfuSYflOqbL/z
E5PLGLBKVzRvecAliOwCP889mM5+6hlTsIXSj7gU0WjrIyURDqpRNZNrMqBe56cJhPZCPOEBkLSi
Wvm/Opqm3NYIX1Y+kF2GCRmwOLZ3nq7+odzPUdAj8iqiyuju90M2QUG97Ryh+oJHG2cvfpqrjRhd
jOIkJHaC1zDolYMP5gZjdFyz3IXKo5SVYXUibo32XMYlmJeN6AG+Qi65KbPSFIK1L+nsMfYo5/Qy
3P7WT7118ye8LPjND4JUUCMTl2Spds0vjHi2mdVJko0h0PAHmKg67BFvn6UOcYpuEA2MPAq5nS7R
C1xaYsI2/8ubkmD7IZp0jsNXxQdgz6fosytiqVf24XrY4mvwwTWz4TDoMEqcgKb6yfwOFDL3CSey
0As4jLl1LwzuAsCN8TMF3oj7k/qlkU+x9/TiJTcBV1cJ92h0cFCAceb+4gteMrxj9MN9deNQEdYM
Xr5CwAkw/4h2m2jtjCbN9RMCi5y/k1pkEffeX3l9xm5ABpICd4oVvoZlFdXS4tv7YNyQuvq7nCNs
CwC5UXEwK32QLWkp1CgFZ8428EZSj3POxG+/9lTx8inXd/UM62GpFEVsOfRheydyRgJQSZe2v2CN
oogaKkLyatn62X5H8rj///vepLaw/aN/Vpfv+eKy3d12/NBNhDrxCKg8d8P8KWRiyOn4UJT+z5Vn
BXhjinO+fS4tb/GPxYh4kKeE1MhuTy2aHTfkR9JlNxfOyavhSXqeo6fGHjBLnkDRDnt5m1XWFZE7
EJQ3S0J97wJ8OogigBSlST3imzgSU2PgvJ1rXobDzd6Q4PNvXsboCaKhQq1LkudKLh/qgz6mQMfe
gPE9wW7WhnFK+ZX0xLsESjdfnPE4z9iX7Gq6zBAmPbqNXtSejWEmVfVoy/C5RMmK43qzvUcItgQY
l4ro+/PewVZpt0ghjRar4NwKvPrtzsFZEdWCVeuIot7e9FFDohPROpe9lbhKVz5wr6dt1ZkxV8tP
1/Zd49NjdAYR9sFXBcKkYMmoohR4FbSgonIQK9P3EmRHCD7+36dGM7cJkMNlV25+iba6u51MBlKq
kcaztcH/djCWs1/PSA3ddFw0UBa32Xe0mBM0jqxW5upkus4jUzwb9ZQzMADzi3QNwx0S+a+SU5/7
aixNFHdAI2nLOH56I1QTCl7slKwkB0JM8b/qoYmS2mdyYEUniawegeDWTMoSQ02yzfIT68oEMa0t
vhJbmV1aekAakVmRj191xWji8eX6YY+wmIsGZ83ajkzRmjK0nx+PaAi4Hv9ZKYGhCfvv+hiqvmC8
HxF/2rOu/tPvswZHzGLixr+v0neP0lcwRl2gOmUcZj1ELi3OdT4FD1MGv/rYkbIrB2skDn075a9l
7P5dQAgGuOX23DDTjL1YADyq7HJwLR9Q9f2UF6SKgsSDj4SjGuBZ0c3zFef1PbgIXGr2ptXC3wTP
1ZCml5rbJQQO+L1EQzxJEBxgX6aLw70y81XXsAR0PEOmAT47aDRPsCf2ckcIwCG4nQdJ17Yqjen5
nw4urxdturawoFeIbEW3qESyAXaf9kxe9dapjzCdcdAGKFcGWd5TNu+aT8KcB6YLbso4sUbpblU9
gb7db3VarMRQpUiz9Izeayn6yZ8z8b21MOfVYCnP6OE/r7ncfLdNyXAJF+jUSc1ltX+RssZdHOSE
GiqcQ7t2Ug7IpRqFOssmQaddFEh8XER5/8o5fFDEj5/j6H/qxDo4AzjswqiK365VzmcYJiCZFtFK
+/bIc3drg90JinuQj8aTf4Uhbob3epv4DgpJOqMxg5GOUDIzwpcjODgsqP4Sq35zGNP06VbgbqzL
uy+n/vR5GWHEBkcVIjpls7FHhs8ANpBGg4zaglUmwabESY3WPi48zqjXl9hQZ3RietRvoeDIo1wZ
FLdJhvLYmSMOL3dKoMg4/BNwKRTpbnh/mk0A9wGDM3hu95Oo5ATPk5JPrk4pMrucLlkXrvQRfUDV
elVsxQqi+ItOQjCuEjh6K8H8/K5ncl2zXGecAZZ4/OFwhm0cIBWEAS3ZP7YBI3xUGXxumVe77JiM
Qi4oMwFYhe7JuRDjbFF68ocqsoJGtKIBTSRTt28vPAOYeosAyAXHBAraTMSaPSkBbNCo8BF0nLR1
pzVLiZ4OcCvqTjFj0QDedwfzVPevNbOONDjHBoqrCK5WstShXxtdPRu+IRIvV5WgcKVQ4FftGeRN
dWM/h8sP/wXWSVLHbjeLcGb6O/0pfYMReqTf2qkOoSnohIutGHeANN/B68o8ZSyZk3CzuQvcqfVP
3Hy36e47bhCclIRwJJmY0ZPCPiPbxPN7siL0jFgFgKIfg+/MLrIBwlY0eJsr5zjRviGWBieQ/5cZ
si8+A4YfgrEhy2uzQ8jzNbPG1YbxKZjVDiVF1dOmMhLytxS3LoPpWmPTQA0J/1m+Tl0D8EShGBN0
PzmRLPMkSFCM2EEiu+3yif4HbK+IiwaMppJg3X4kDbnxSZdijZb99D76I/TseiPQTklYiV3rAMo3
M9bIF4fYJygpJaSht1otMoYLiA0z2+y40mC5vLYQIwOImuZPXKmIPkHn7w1WjJax7kHKG4kGsSBg
YifwqoRCXcxO9V774Ln1dANGqtNSIApJYDzw3rmbiotBnoWcCzJt8HP2QN5nC+rmn6V0gGc1E0RS
hRBFi7pmBEUm+TF7APOLxCmhSISc3Na4/A0VtXPOdq1K1ZgmjqivTjhUmQNVi4xNDdbw8IZ/fwZe
a9C00AnRbOGGytq0FQWCqTFDHgFfW0CnLalpDQqrfeJxAif8/NasAmb+XbJJP8T1xw+HXvdHYZCn
/b7sOA46nuGqmt0e+Wvd8vmJt4umlTXmDNMMkCnhDhDymLX3JugNLBOlyOpJALqMbHkdBDplxgNC
5+ifs0Y3VLW7DmsXZd2WusQ3IdhLoT3rkiUtcCFiiLIUjD2ZnKSrQ7uCN8kAmuVa5HRht1Jize1y
WAthv1SiQxMXdaa1WcSKckB6LxKWebjShaweku35U/v0B95HZAV0xN+ANAeLAyNzPKPRIF3gh2Ve
TcYhA+O46g55eTOugCUrgUYQ+K0mpYxa531FEb0iiYaJ32TYKvqI8s4ZPSU/t2LglWc81Wwhe3vx
V2GVqX4h9f2m1KWPe888ZVXQ6txxV3lGzuaaa5m7GxCTFuslW8iajYOpNcL4ZfcNkphFPWXezyEL
PEimobVmVU33I8lYKMH5QIHHZ+8xAsUO8AK3fESopGgJIyCU1/JICpwUv7yrgIURPdpqsFsbtg99
fvS2pIXtB11ju9wWau0jJeC+iglK2FhR/AoumtYbH19J4YA4T4UVGt3sqGL0wh+ufUuY5VRc8nv9
0vKsSD8XpU+ycGhUfQk5hKz1QnssYB1O2YazIZDBYux561zOBXlo+sSh4vUfcQ9x5wFbnx2Eg7q3
ZP2qli1QAVvwCpJTdMZ7YzlSXJSAFAiqO1bGfKy8AhZQAGdy8FLaJUPPACexB++YWwMJrwjPvIX9
ALTTuX4pfwJw769aai3fMPM38RBVBb11CBVhkgfL50F5pggysXm0hCKzsk1aV1WRFkn7Re6+vDDU
BwbllnzbQUIsiKwZwbF+/4Up4XMsd+yMV8Z6kdsiHa11Azvj14c0HokP18WIbHvFIrJoQrO1jm7i
v+mVFoFMgkTjxExt03WY+SGUzIA7NEid+Jp7fnGXtuFH70wKIRjSof1aTo7j5TBMaf9pbfYLQAWj
nwfVgtzMt31KzrswYimbWZQSFmssNJJkeOl33UNzmDXQbv7qVkKYFM2ZaGGVWY6P79WrumcjnmSw
rIJ2BKkt1Ax2bl6cDJz2qp4FNdNhxznGQIW0M1s16zPFGK8tDbTwfxR1mswC0xzbSJmdeTaXTcRo
ZndIkX0nKWUvconqykYxBkn9j2If9Ng1ncLxUAd/Pbgt3+SIxLc3pQjOyeE0u3D/PWmozU27aOIv
01y8VVbahcKoVpcSU0F2vck6yEKlIuyPkXQsjR9yWoGLZMnzy6jUnb2URF2bsl/Bhyd0Sa4t20wS
WCbElk0SaE/BBvgjiGAoNXtrzOVMBXbRgaAHIbftCeH9q+JGv6MeDixUl20kpWW+lk5t6EjL4ZaI
tzArPMEDS155mrdLgLtv75qWC5Y7/TeIucXCZbU+t/xbU+9+ZF+BbaYjt4yB5T/OMcxcLzHQX7li
4xmAoFmFgTomocKUDgykA6ED/FTqzZwqg5DYRXPP7VSNfOazsOd7kKtyLT6s6Qzo0tJRCqOqSVgA
kqv/ndqTO/j+TUttb6RaLAZF4odMhnI4nBeAnwNCwZ0GOatdPE/AC8Y/JrIHuu/POeVE6A140dWg
CQCrqV5Fc9z+1gBVX0Zh2lulfHWC/aOysoN90Ll2Xzsqvs35lnSOli/UuBUKaB3cAjdCd8UERoEn
4C/y+gwQTGM2Mzspl/9cI15vCBKfj7F7yttZ76d37jhP+vi5jNns6wyRwR7nm7E18P9q3rzgFhAo
tjkZ728fa8+fSpZ2IDG2fXt6LUGF+LigpLvY1eCvoNPIbKJB0/E0sKCp0/mQiyYxGGz+W2Zt3yxM
QfFqbClV+R1JwkhoMUJfEoamL7Fhi6u9KPPP40fDVMRZ6O9Vdu3R84HqtVnQ9NlmZx8U0SWOiIJq
5ykI/rEWW1D29L4jtndbcaJO21fPO2gNDynYD5mvMTw203GPAR/rN8i0SK2rd6LZMBmZQ2Va2XOW
D6HyuY0cpdO+MnbUVkRkfb8amSgx4PRiBOZLgMJTYosGUjDOOF0bqcaX41mQjKIZqOev9+rcMWCV
lsdAcNqNhrkzkf1pr0WoZvoXsh5BHjIFQ737JZu+huXrDdiQVkYMRPyZ+sbRMREw0itSW/uv5hKH
aDvDNLAD5nntbMlnuNF1yLBG/tIBcGzhnbtQ0Z15D3izfgPTcQkNG+FSBOFxVG/oASgJyFdN6RDi
ckuGH1ETspEF4cTIRzubkn88Ei4DTr4Mheo+sCHWuc/LSY61jY31oDX4pxIfZN/EpWm1zu3LSq+o
cWzlRPwky0b0iIRnmNgYrOYcKt7BM9OLXi3VBKkgDp2AAqMTM6XeiHK3tzOyWPbwgVKgbUWHZSrK
WzDGJs1pZFsIIZpGJiuZFjEtWcnLasPag7fEHNjGEKkfKla/wXhKTIRCu/21csVhwWChUSaLE1B7
8qgl3s+fD2yZ4u8ly+mXXglGpI6PQ77Ia+CveUUrpuEWwCauoOGdIoIDTBzFiVstHuF8/vwm6Lqc
kvqtDvuZgn6orFKyMGg83w9535ajvmpQ3eGAHBl39ETpyeS9+G2g4QsUgfln7wWJ0Wmwro5MiHb9
vvDjCsBqEeDMKjPI4bQYwr0mTk/Bn372ye6ZyswPugyEmpJrlqSXfm7/JCoQytH1PzNn8YY56PLQ
kTbVg5BHmtz/TEq02tS5QTpBEiGNQXXUkAUw4q5Aokddeq1+gesP1AoyhSqj/6V9pXl+zW5N++cU
kxeySto8H6dUJ/EFSwuOjnyXNvU4RHtp1AlPrkz81W8rGIHixYVlodb1SqzHmXgdJTX7tSPJYVlB
FA5bJi8Kd6nBsgISlJxWHObxgB2pL4Nu1lthBumYJlAblybUg6sFhcRQgJAY5O5ZBdrcGlxuug8C
ALxE8d3FbRJOx8+HgsD2wsQ8fOIZrEanJd6fHH/9c/s8X4YYQaXJ15a8FxiH3zI3XAHwAG4f2orN
u7rVTdAV3LWRHJ65HRSqj9rwi+Ex8tZfGm3hH+HRf+HnEOeeaUuwktX1OCTE6LjPnzWs+u8uKMra
i5iQy7eNEY0qwHtykZSHnmb9UBtqefRGEo+5H58onqPT5WUdc90CgOTqHDNLcEbJGCjO9PmyOh84
8CPdbTfjH2lBrG+ftynMtghpu97vDxm2BKFXqW9zH4EkCfUey52YfXVM+VMfjDiN3eAgbWsObLUa
3j6GKeY0WzKXXvMsgTnA9hI3bahIZGSkL9n1FKHjkU9JvFuymT5YZxEMwuQ8MZx13lejOcYpXZGd
zr15kapW7AUAuzfW+sbkUZJLQYxpu1szBbB7azPHu18G3eZK583p1MQQxywZ9PRYpvuKuHviU+e1
tnZ01gNxzvxjcKXOxG5P3WLA53YWCMdmmBSqKeogksSTY+afFd/YddN5L4qFdF4mgVQw1Pb7xKo2
t19pot7N7BdBw6YzYHFoYDKG4OXsESSt+IQ6QF+F3HLj6TLvcI0L4L+T2Rsf8Pv8882sJc6P+yti
Go9YNr9Gkd+O3rEa9C9Z7fQMU1mx8keSiLSJHjyN7j3lnv05DVEHQtIX4N29h7qaCkzDZ9ETrCI3
1YrRBA30O7GKO5b16PN6/CRStNjHmddQRUetM5XAQ7O4NFdCFwjpB7cs0uP+1lUusFN4v7NkN2Jp
dr+BHY+1qo1+4ggEPDuxuN5jSahTERHMTOLHnkOfjvkroL0zq7AxCDi5V4Wl6idjMuUmtMdziB6J
ir+rEFG+qUqIB3QcTsNYVDLhMrCMz2mm9tO/EPdUWI8+08XJ6Q8fdavAkrTPMI0UzAyQAogR0/sX
D3lbisiqdaqB5f/tjwN8Yzx5fPvWD381vlHXoArb2DjwBNK3RAfWNZ6x/dJIKaQR0fj4fzZpo0V/
J2Iet7pDmUSCw1lzD9AfEfJ1NiqVQ7XHKvfv47gxhE9YcDKMh2Tg4XK7yTfqnIP4Fybb905GXLDk
XE7ev6kqB70V4vsDzklJosbQm6KXFECAaMbJ5nkyWT9AfYZSXBJHMq456AU8R9X8iMhoSo0FlszQ
OSWyi+5Fzh1l8XDYIiziPVC0OqDCsrzpW9aUaQJj+F3h4XZARdZ1iwkbkszOgP6wbix0fAjpJJSE
VaGhbd1exqHvAvLD31/w/AVNkmxivwqWJq/6Xb34AahFV6JF0EYDqo90EcjmwRT1oRjSRlLq4rU3
JKjRT7/x3zb9zDa3RgOT9ydSd8BlWPian50zadJl+BylZWMpOtZc7Q+0cRWcoruPAefOO7PZ1FX6
nUdyZx8V2Dwmw2fqsLz532MvtvR7lyi+pxqtQmqiSPGEPN68fBzJkt5TzmeDB6cGtsN+eQ/evIG1
f4vpC2R5Yn0jKE2HVbBbcRZFor8ULm4+omZTkBkRMHVCIQ0wEaEVId3tqrotg15MlI3wqRkclXpf
UUgVjUYb9p1gw7c1Xam5u5ll3nbWME9d+zNzNlQsoZ2QPQi+Q5cGVgQcfnIOPQvYPEqynRNUJTIF
bLph2cTDQrsTUstwvFqClDACuS8AmIcGwh9SrsKqsXKT/XuoVAhLKqSAoBcnprvPSR9uqTuljhwM
usmZCuPxiXZdZm8I9X2OJufqbWdZ4Ej0LkO90EdmV0ixBr4lDNLIpagdLpslFxDOklM+sUgZa/fT
1qEqzR3R67QDu2iS2PG+FspWB09zWe2mk6SebMI6LTf0BT+bv1dXjVZyHy0+xU4zfmGktdmmzUro
ud5wqqzinwnF7611rd5t9O0dQflxEJhjKBY/4bQ6fAfQL0pfYobxED0z30t711t9v/1gHOHaT8ek
gEmPSIIsp3qhxjrkcbP4hCLmmpBPYLvFjfvBFgKmnYTz9+ObDfH8PoHIckzjmCXBUizYPwp8akl8
r4ZEZUREf4BOkpd9OqoncSoRuJWd9e+TbUucIC2+kW1tb6Ukn7t6Sykw4clr36XhnG2bYrMi1OQd
tDNSJnxRcPPXoq59CSXMj9RIRd/WeyUE+AaU9tJlgNKkJGFKOCxsg4HCe29wfCcSdbdy3m5zaDpp
iYwvv+HErAwd7033DhKDGMSxw3FVX8XqM26qcChDiC1r10jbpHNLXazBlH8x5SlE2qnfLbgCXEAU
oaXI3nxR4qMI0RwafETqU0xrrSzhgIl+EhqrvnsMgLmn+hU4ggp21E4yBVTNTTTrYTfw6HEkK10B
hFR7J/Vl0CitCeYtyYDmHLhxIQjev+mmrctVeVfLTuur4dEG74EhY2KmbZY6E9FHO1JGkyFqRHd4
aiHHEISyJetGbikN893g0gpw78AWVGe6eb3PnrGs4Z+khfdD3F2nZlo/3/mkpXcfDwnVf+m/n630
GdFdHIgNY3/g4xNWUM2zp8MIq9zayzIdDKsXgWRs8Fe2oY4rEiL9jKh3H4PsoXbx1Q9dBvDDemo3
MMzw/2/iljXVw6C4cmEplwtTGxcpXkDhDMKNZnSBkoSu/uhU7xRNC6nJrINyP2p8eFctmMWLBODm
+GwzYMehz1bxUpQu4iJC4daRhIPqATpqtnU9R2O8tugbD6eiSl1bOwUu/N8vn+aXOeIW/eQuVZvk
M41GoKX5w3YWnipev+AwUmA0gl4ng7/CUGfyAzAYsQ9swJakPieCYrZ5KP/YNWbLp6HP6bejYaVM
DJMa+Zp0rHPw1WwJ7UWl3XL7VudfNnh6MDqGR+5Aq3hloM/srWAaxfYqXuHXsmbcu/ORc99ny3w9
o/2aFQGF9v1+n9ztLZ90ynsaNquHsZRxH+dv+J7V0kpCGP05Qax913OrNXABTYwS+/TNGaaAcKH1
w4pLX0CwmoCIVC/goMKVdWv7kbC+OL6152gIJ6PWTUG11o6T/ya5JV0dODn2pkZxgHETj76qN0g5
elfX9vMmjvys2JMSwRF884f5gt3nIPpkN1elZs8au+LKCz7X4VNr3Rsp3SL4J3l2IaCOP/uM9RGx
KxSZmLIkj6EUSY66MDCQsjfT3N1nom2nreL2uLhrtLiKJuvtdjnBQ/EXux5UQp3AnSNqkj4m5gXn
omdJjx4gDO1KYpXp9itMhG4dbbDKvFK2FJhzEkWPJNL5sO8lJZyXEzY1Xmj00kiTQNqZ2qTAFKlw
LPOVf3UjyTVyaBd575L52aM2z0plXtzq4CS5G9hA88fyrSLuYKqgnswvR0xMxpUcL5LY5pEADWIL
1p+XS18FZa3oYs1dNxWn1pa8Gk1gItNUWUo0ojz3y8RR+mPXNbhT95E5id8rU1BAW2ul4a5WOMMS
Da1c1opue29gEOdIFh82rQbrvdQnRBRyUvwN74yl3py+Qne7MuyzrERz9HNWT2yB2vRPGcLKjBc1
SsoYe9VeQB8BiJAY8FTNB9NIfUNIup0pVYc7O5nS8/Ed6sGF6U5DphBckQOJ3ZsjWru3kJEqbDg0
UDQIbbs1wecUzhhCitxsRt+w8D0lAGjCs5PiioHL+4C63p1OSh1HcUD9aXzw3grHWagMSWYxeDbX
iSwlia1bQ7J10Cs3vKJdXreF/PCsL2QPPA4LlhS9WfwWQk0ucSZdAE5pWQnYKclMKDeGT56Tcs6J
SnVexJHGJOZ0KfYABeMcRxrzfttG9E1ruuwe1h0OezdHUOOsVUAXJ4gIOHpY8+Q2bH2TKBrAAf3E
49bSsU0SzmNBF0f2nUMhwDXp+KClL2fuh+Ht/po58LiKix7zvkuW0p2J4MD5604AmIXr9Yr3qZwP
cPGC/T/ioNfEGm4/iibIPDOxv0v9WBd0+yUvv31sAMZS6cGjkd23ANkwEQEaVUsohQ7yD48q2sny
D0mVEbOEl9qA1OQXmFHmNbD8cZMz72CaBfBazvLRBibqMVH7xblSuczo50RchwoXjKh5ApunL+pz
hK3+kZFZlyXNVEOcp4cxSfZx3gsSb00/PBNevsIsg3ZSPCq5WBYH5ryrjZcI0hAyaUoFpqw1ks9H
n4IX+Beh5IDpG77YiUP0tW6l/h9bzGC9mBtr/ydSurGvLRdljend35U3D2mPSQAlE4xhqu4Fir5b
kUcRIlX4Zvpp5niyrG/148uVbIEY9mqL2HGCI99qkQqTqkk/sJifmeALa592wy73v+9/WWzj/J2E
VuSAmEunPnccEbdP+DK/QOpWuvnZKWIvwmFEHK718AGbkAi4n24ZIP1GvwHDs6eH20TtbFZ9PDDN
Ly3Pu9n87NnHqMXa8wE+xFP3izfWOJo8nfIGWkz/D3+Ct28FdlTYMD1gCo4Wbpfplm4B2Bi2HPht
cUZCWzOJBBvqHvGZ9mO4s04T7xPNmQRV00qcg+DQiKb3g0/JvQl/22n++WGIvnhJhMQN3NJnY3sv
4Z/bDCSouwszuQz3kSkTylCnuPdHciFcvVm5t04DDc0nQcPTQGZkqtiVXQEMuEk7QzNyL1eL3t0U
CfI/alzmV85uW758ypTWSIstGBzcyzzyghUuqLjaZMZ0RqmHBuS12Imk4Ir+ispc7wIu6WYIcqRu
+dgcje37/UgNABMSHqsuIJGw0cdaPk7kwPCgpSQG5bg5zO0VLXR38QbW6h0+6iQCJMGnVBXlzx3Q
WoN/6yE8KPJ+5uTZZKm+766RbfFOzy2FgRusYY24EdNfBynhCllaVkhaXTreQLVEXSkpT0MY6pxx
9n6fkMo6EuUT5kOrFQhrTO0IWDoLcwstRNl5u8knzUPfNdZOxC6h8TzTWy3wP9xIdnDZO1eclMqd
BbauHWzijGTjBwXYutSMiNvSNs0KZFihrYwW1gSjQRFVK0IW00hhcGUJf2+qqtUdIU83u+M5cNfg
EQYzxElIom0Yb7qYwZY3iENeVV3LyGNHaZnGgWP77NG6KQ4x9n7CE5wbhnGEKGzspNxXM8mToh+3
kOmfH9o32ZQz3zagXjNr6IE9etpMGrf9xVwxegG3nLRdE+M7LSfarM7UYmrrmlKUEReW93FVdoaa
F0khM7z6vZ9jzOdyYk0dHWjcv8nJfHkQQKbZ39r3Coo6iZA7CdiF4D6sHYLorz7EynJxwQnyUvbG
NfX1f+2qxrAp4yJe7nWR8A1Bc7VftfgaQ/je3GVskN4I1vRa1V5EPAw1pkwm/U4HIWRWuUNkWZZW
uRQ7MKXV5aM5tHSSbpwgPdEiseZZNKECnAWNkgFgoYhaCpc+7jJ4RWMJrxDOlSJzB86X6e+SVlLU
LhKXxAq1B0kqVRv2Sb0cuLW66y6U5arlLGSzd1NR75qaMF8lsA58Y7NeaqRTe5rBgXqB1Vryn/DU
48f5J2phohA0CMx0zD5ZOKRt+28Us30/wuAzBG3RyMpj2DvD9k0AQ4Fecw/rD7v4aC49o5D8FkC4
WzTCgGCCHrlZE/0v5h/TEdwxFs2yEAgUf5nEIkkiHIPEdJNqnAjkvJTCH4OAUDJT459M3wBZxANn
T7mvtN+TQst3xncdh2ai5D2ugJ5RpQ0SLJnRa58Ize+dJthvgcMaDBEe3f65dqZtcxIJQ2qN6+Ce
tzcUsUbq53EPuTrQ6PmpFF0Wcb+soFfRhpCvQcdlybZgZ2XwnI13vUZbPZJZeA4yFZPjyTOBponA
ngN5YHTo4zkDip/zZ1s9SBkYI0OpHw0x0fAURPOg9UZOjHs77mmPhh24ge6AXLLHcvp3HtkA04ur
YoSElgtFvD0dZyIDUOqt4VF24j7bfORyT6mB/yCvxbIGJTa6ygO8dR9esvXmrcGW7WyKKO9zcoM1
jyyPBmBAEsA8TbxwsNeq4XvNC3ogThUJU2tGVbOFHfzcVKbEJkKuISU+ED1ZOUYGNGVBDTFhWHm8
pxre1ZNpR8bNDARLr0ip8XtM0Z9knwT3K5DJGj/diRWgRUmj8tjGs+ORyBQ6XOnhi4mD1WnH+Fw3
ZS7CgrAmg5JT4W+xk2D/ZiHOIGdjB3suD91gdh6tp83Dd79UiiNPLdAkNBks1kFy8b1fU/CwR1S4
U/5GSR4hKfKT8Qqc1dukT/F2czIL2Y5Ly6LMg6bOp+w0MFqKjc+5JCyg+/gzC070eutUjq6HmRgp
uVxdALsHwdWtV/Cy0eWSlrLM/f245LbImGPyDwYkWdTIb+b8aBjQJ+YB0ZHo1Ddh8aqd9PVYVgEr
IP6sqX9JP4quNfbXj1OB2uQ3/SPG4hLC4lDl+AgpEw9zpMh0tKGg2B/tiLZ4XkNNaaO3G51r9c3+
gE/gnn02NMbAZZ5CxypSH53+j1WZt/WYudws/bQE6ry+hklVsQkkZdb6T+iQjq7iy/EYJDeejwba
1Uqnpv0xWhLAJi3v0uDI9xo1nNYAeV1cRsPQM8hPXqLbjgsgsPtrgF4TNr/zdWS/emoNkZ6ZB/nr
U1aED6/mYkzr7KtmXGWnDWdy70e6Zs/JgFSeiNT7uxoJ4J59wVW8MiIpPTBzxbauInyUIZiF92sY
QMqhTryEUsmYmJDjdYIivMRPJHtoGe3KMfZzvojEuHOuqrPU5RRN5eWoccjetBVqqMWeoC2Uzvej
68gWdGwj6iFbjfqlqCq2gXWrxK/FlrcVV6uEU90kNTdc+N4CF47TUtpduW6BokDhsv4np1knqVd3
LJPNwIyYOJ/FiFYcpW+k55ISzKMakS+8ku7jbknhVDaYOX4S638ARDJ0c7zGy+EQTXhPZmxzP5lo
bFXu2Ul91O64T5L5O69Zv0HaXBgo/ecPU5bE4wZES88Wxs2P4MSaVHfK3uDLsa4xTj11+CgxFZrQ
UkQJVhnB0poMqvOsorVLw1NhBMuEbhZdo85s3Ty5I3fehITBJYZqD3ShN9ZZ0Aam8xEb/3S0GLjM
YRe7kDH3eOrYUMOc6mmvs9360QbJ+7XWOSuDLHWslc1ONAaqqbygftp7ZZobnK8HuboUmJJIwV80
iBvvB+wDEBvo3f2jq/3eD4OAcIJXkvgw1XNWlzFKeGnO/cqfZlhlcx9uHa/rgXBD/0vC9/xi1YaR
KQQuUOvTUcdSCEz8bsqxJYw6EKzu5uS8cbcHngBCwhbelZoaH0wkvwUc9KMTEaD0SCC80uPuYJGi
LhHeKdEiQm9NzqME9eSml3aICHrtCH4c5ewVWZUhMIQGXUMb5T1ED+htL3yTUTH1M7DZ0MxKSXa4
9dPWHsQeNUViblZ+m3zyUGGvQauvKwISsP520YD6JueJnDqYv0R/hkKxBwNZUCb++kq0xwQ3hVEF
HU7fgiACKIs+y3ETV16XmfwB0/DtT0yUKqF2IrhpfVD1ihqmfdZpOVJoAS4Wsj6lorePIvvgio+o
KP/Gd/ONxFwye1CtVIHH/lyG8fdwbI9bIsNdMcFTl4DKSuoMh5ko4XZCPFFSFU1tjL5ewwuU4Gff
vaUUz32H1DNcbsim8Vf+ZjqbsyPpd+PHuiwu6pXJr3VWYXkmD0KtHtEgkU6qnc2hl1KCQpT6dCQN
PvvGXbkYBk9voAjYOEJFStojJkwor0F5HvkJq+6e+rEVpIYbiJh4Vzk6DPh5xnrhHQfW2Yz96V3s
rk5QwBCvuL9J62X453FmiUvORWyQ+s/N6X+0+6ZI0Dz176luu85oliellrRAwfpv/ZpUWTBFCAaw
SnQ27qKsqb4kb+oSwqQoQ41zaDMorKXINzc0Dpv8MXIGe1ST8ugO/jPy/Fg7jE+Rz2VmOa88n0Ee
uH/82kvekKSWNX2E2HWJeWrIIWz/9XVBxKu++3Ocpp03wWDVBxKfNPizyafM9rxO0m/sdF9rW3Xi
o1LA9eEQL2Rfct9G3vf6S/+x7kc1nrklzLTeGhD4OzHMBzbyUuTg4d4MmhkHp6G4JqijpxLpm7hH
RygJP7jpNjJB0tRcj29Lap4qOPCxNr8zSfREiuknxEFK6DcDBOlpush9IJGN7sGrhaI/G5OiBEHL
wZkwX9oToTJw9+FGUd9hA3tHICwNd+FVPIYMcep11warmtEHFXk56xmIuMtlmJapgvKFg0Y5WP97
IvKyotRjlcPjph6pRtxy/+x5/mA27oOsAFU7opsJHd4AzmWH4fZJI5QAtrn6RSpGZpqJC466Djk2
/tikNTk73GlLMPslpbNZz4iwypJ84iNVmJWNCO44WSW0HuHkLNY0AY9TcTL+m/JwEKL4nBCps7nu
+EMceyL5Cd+mvrI76VBp430xm2g5bcWAI++52EcJU+KDUfK3DwhdG8uCYwWYWaamN7U6+PdRSGMG
r8+osVUjxxzszZCMN++CdQoc810KubHhKFn8Hb5wDWtWfkuA0tGV1C1XzgRApk7Oi3hdnPyAM59V
Y9/+8HlsSNb6g5VOziIeAMcKglahPCIuWS5OyBee0ypAGTQR9MNnSeXmyomjJJTCVDKmBSo/1s4x
w1RN5nQ8y8mR2Uwb8Glk5mAu5w2O/8YnACBM1F+/v0KTYnzyWks1+AFKvVzXgTcqtfmjG7J3DELi
25sjsu99Z2rwFG813flqlhwfnF7BC16j86w760aHgkeogO41ESd5Dcx2LS5C7p+f8/KvhztWLiYi
BwUok9fORnlLGUohjoMx69L+UatgOb0bgpXY7JKwf+PY86cpNrMusEvPYPobjRYONRjwR2SWUubw
bYDNCVCADPAIatgPAEXZUdDMfMa2w1oLi3K8yMqNrDR059A+q6utXAoAzypL5ECKc+mFDXlXzTDG
RMCtCwEpaRtWidriyi2HLJwqKwS+F+JVgTl4xhOo0pAcrvyNVLv6We3cZ/+nXrBQHnpt5Fbgp9B4
6Q92o7JZz77gXRxyTl0cbmf7X+49tONhM6MGTPmiUrXfBF/jnv5Omc2/M4K+V1bFIu9yTivomqw4
fdfdG42io7P0XAsNaVJTs5xyuUG7HkLleMY2C2g3GtHGxIj1APLUgSeyTJ08LpdYZXrkvRGuR8lm
FYtrao0/Swa+315Vuw48B9/iUp/vme8aGKNHWEIoh+aa9SPNE8M77Q3CjQ7FhZ5RSXwTAesj4g/h
y2EZh/UnwClEtcm7qKtEV8+D2F9SBstbheHFIOAsgSkXiGTmhTlsaz8ZUYiNXvyVnlFLZdxIJ3Nx
BGPM+ZgA8VST5U/MI4fcjj25n/VnPF61+6qFvoXVvIC1fmVJXE7Oep0id7lcTpquoZJwpsPV7kXR
P/K8lgLRuKFQKAziquRSvmv3Iq1qQuukIBdKkqjRT161Ww2bJasde9qG2/WKJ/dvlFTbxt/cuFke
Lyls+uGysvfPHmzqLn9AhMM7JcC0CPMEbAg7A+cGmPPijfVH7yR8AEJ2LRqEUWVZP4ag9qOoEwkS
8igNHqxejumLzNLaZEQgnIImSpb+J7ZPHr0IKsua7GPjcuKVM6o7w48Bxvh6edHGumeLTi3+s/Zt
lo4xQ8zp/yEPm/LHpCXlYJalrvnfsueDcajNK5IRMP/EffshfHi9wXFEHAHAaE9yqkDvChmvkUI7
DcdyBaUPdKFCaRSb/So1WP0GNh1IbWaOpkZonGZBzSHIClafDMu7Tkk2HfMaMhF3WoMsXGakNe/y
ww5C6SmViR6N/DJEOsvtwwX3JtU8kPCFtZA9Ka4PrDHMSC8epZTUtKlRDHd6FRz1G4aQ85CoZQSP
cvNis9L9GbOtunXrbo2E9hpGu14MhSPqiCmCQfnVATLwM2+L6jgR5/nDou0a8uOWdBvqORcwLbOI
tujWtUpZ5gcrlLxa9zdXG0VPWwM3x3HOsUZS8eeZ+8qSb07mZRQcBS+prIPVyb1d7EPywv/UrWwd
M/eXg2W5YT9b7XHMqQsyXdPcQbzdh7pSr30i1b/pumgW31PDwIrbzuSnhVY1wk4QSdvlySPENnIT
KpV7EwhzJ6rgoZ8eTWsaQn3QkKWBnfIVLm9JQu5U3SQIKfxNWY4ZemexTVyX0GOF3soPboS7eS+g
N0xOgzGNcRBhShH1JnWVJOtesB2holBV+OKpvPdvUFKl0jURKx/F4cA+JeiX8yp9bFpAXe4IKWUg
IlHjPOGHodIwkRM0ZQ6RSYY2/uBAyjkqMt1v0kBpu4kYn58R/g8ppOD/QcsaDSTXaagJuA90ubm9
SdERGdX+qh6SWLXBGh+bdjEzMiacrR7cdr19ZEqhtsPT2fFa5ry3op1Wh+394TJcaxtLYg4Xq5tg
5Vj/oasCg92FnTqxCxUhNtHZYXQK2is4+KA548/nuCZNyT+ykt9etvXOfAIG7oEfEWEjdJyESzX8
34hdlhHtnn6KL0CXCgJs8qPyZVplSV97JfgjYpZ8VZUbXSiOiUj+hrUDluNiUiR71I0m98pKm/MK
+d/wutjzIRgxG4ZgmU0wDe2aeH8vWEQhjxvAmxyuuURCnLWqCULXXaesoA1Bh9CnpoNyoaraNEID
8JrLwb4ZhSvOY/dqkM2GFpkHySTUWQRv0Ep3EI9RCps9PQYH7E6FhBodqtyvSxc6HM9wARknj4uh
kd7B9rTNiI5H8kDPYaDiwZDWubacBh6AgCf0rVfMDb1oJOU6ELCZYj6svnEFT7A4jDPKhiMdDey7
TcX8pCdoL3ali5zKX4pdoyze8UhARq1ALdW19oC1nOgqc/fSQmmq2doaOw6ZipVW26oM/LCvdXyL
d5PAjtOZgl+NC01NxGjUjbQ7O2lXDtcYN/mRDGZi6o4+7sGWPt46RxPHJsl3954qfE+ayS9KGXdb
+2QoPO8VNRMoZ5qrYfujOvdSRUG2x+pTE2/WD//woDZeuboHuyCArW3JHyCsUqrrUEDKF10RRGJX
gARg+bAFbbujcLMYNr5RhcBbz+eLOFc4REaiTOC63eELA6Q2+J9LiUh9P3hXnYx5mpBsN60hJa9N
fKMF8ZOMZRckwdIZBsPWtch3mdgrg7wNmVXXD0b9dIVYP12TI8QicLaq6sM2ZNQidiOV0Ynb3i94
dakDMYtXMo681TISprTkKD91FL1ZtCQgfkIlwRvhG2Jxd3MPKROp4EQo7w449AuyCDfNsGSdWxvB
dNuP/lLTRgv3V/Vtg3bdw6AA0ZLxq8AmgdLCrRPKv98t8Bp8MS04vrgN++mbOq2P9mwey+NuwuzF
FEPnmDs2ava0+JFYpWf4lBjqkWO1yqL9lxW9knj0RivZkXJuNfJ05f7oaH39huvPub5cHbJrpH2T
gYgq6UZSNjhC5rZU0pOopLqLhrUEWR7CohdLwBFL2e7c+YriX+nqdwsgXq1Ik9FC8Zexb8Jd1oZu
NAqOjtovlPUsFODhes62+8ohDwYh9beBxXRuOFQX/QlOf++3EUPpibe0uy3WCPSG3Tggckmo9y6V
ojVTmiCMxacFvXmDcIoNiN7nAgD8AZf0hJ/g4QurZV0mwK61Q5u9xEYYTGh4ft6w4MbejN8Mqc2i
+Cf4W/bafiqcxc4kXrghFO4TnsYO93rt3hTK9/NYISwGPZKSrbWKwNcOlhWxl7+loNpcFznN82Wa
6jwgDQkC/2bLTIveesjX6nlCC8S/owaA8kQrzRxUHmYR4P4FZWKaStVbWiytHRGjAjIveb3kXO1i
5wt94nmGvaDjhlO4uUFN321k2AXIucquSWQaUf/96uFIA3v7gY8g7IRTaT+rhQxdnyAjYdtYImLT
A3qLIztZ9NXrBCfd1EBjZclkgnZgSSYformZ8z+/9mfX7JIM08K5MzUE8aFEkveM/CAn0ukMlw/I
2V6HvXObYCVAx1Y64ukGnTFENJemK/wGGSuFOCWR2ABT7d5iwzKGFQ3gQW/SauBaKGOGIQKxu7CY
na4urhT5fGwjiL/Ivwn1TmP6J2xBxDfkZfbANB7kxOEuqvg0oBknDAoX0X2yM6X2mZfMBiUzGY55
0x3TpkUPcvIvyvSdEH9Z6VTuXsQL5339p9cLovvUuQBr74gG0uT6a50Vt+bay4Kz8SHCn4TiYoWM
RpgHFg3NnZXK7/HblyC2Cdsb95T5udggRUoUMNK4+Y0EEHob9SuWoWVOMd8ZEVsl6ZSNB0oMuTLs
BTPquvXL0eaezUwbHBhzr9JNz6AntHu8OU22VciOrEPjfNRPQr5UB1U6btBr+9UiuduXBNrue1wM
CNqf0T1wDX9hZ9E/F5VFkcTawGmh6LPBMiYMSGBlJR7Q+Irr9kYLQ+GPIgivH08k3d4xf6Ld93Y6
YVIs9k43aU1jAmZST5qOOu61pcE+nkeARdtnqRmxTZ0C9Ml/7YpR2822APhWvTOrsHXOEXdh4kzd
Bv1MpQ0d1hmS3GEO2mge2goCZd6hXsEpB7J6GGTiIaX7vvTmlu1/1Le0ZLeGnOl5fFpFBWUzbGbt
3bm11YiCIw6FwbiMiZ0OHeSx+QhC4TcMRej2xZQplVtwF+BME8e/PVMx3mDLqVM1BYBF7K1fAZcT
dzp6lwHfnYyMvWxm259ftkq4M8oxK2TdzNBb3+fhb4p8UpCHs3spF1HYQdhXdLPkCah9imrIOCDE
clKLaNRfinrfb6ksTwnTc52NSxIGMFxFHWPO1nyqdTF0De4vKOb/jdqqS//reoI56CsAsZSU9ead
xAYWMMTtbgGwMGdb6sGLozMMVSFHRJEBHGxwgJ9+9mPj5QwQcQrYFpWkvO9F04gcG8JhCK+w/P8i
qtjYrC7GoIhSkBC8ztxrR5NTqN1xPUWSq8gP2l2YHWhohT9/xamxwMV2LkRZmoqB/RcS2/ys/yZL
O7KKPzbycY0JQU/xOb2OKjHjv5tpXe3Oh6q46RGVN+1bzrkwvVK4jALcI/hs9J4W0lnNHp25tCAQ
SexmmheVNxmVMVXmGmipOzui6KKaVNC1DTGg2aoOC7DkGVmLeZWlOATEKFzp9C+kWJhFO6odTByH
DQq02paQSugLh7BjoJkmvQNSiXr+Le+OdplezTLPhU5F4bD2fprV4GcnkUCB6CvAbh0rTA6uHM6h
thUkIQnS5unf5QQWEGZnYaALW0/6e26inDrUUnTV6NPthPTX8ITHxPWDMmmKNIp6AJSCFydOZtJI
39AKquOGLUNPi+27t2snde8OwdJsqzamE/7Epgd8nX7lIc1lDFYYGMkDZFtG6YmczM9jBkDtda7M
36NcyYMDLXfQRhVCCFlwDWAilGikrw7I7A9ZA08BNvNlky5dNKA3JTWywQSfS3qJRdkDZfhduAlw
6GuB/BG3K8vYmRSdeE7KvXAbwroxNVx8LF2YesdRp5S8OqcK+18PwmPWEqas3PUQMF7pRN8t6C6w
2/VC69RipmdEkprcvTvuCuw61a3AEEOiIAzvMozK3IX97RYTdc2Og8Cj3leRqecr9UQLAXokLWvM
/GRjtfFm3QxuqRb0naaueFEy1jwqtQdiJrTY6zVPGGG/D8Y8rcShiUcLbi2CgSJjLTYycd8i7QAr
YPD6z12pulOS3ILmbD4RXAnc/PBtP7Jg7ArDUCBGPzCwhLE76JKLSOg20SsEBXKAketE6Zmh6ZyC
YlYm2TwvZc0rjkB1nL3oHyJgMOusL/bjeYw0aE18qo4GJTBA1Xv7jCRwboWW1YuEZfxtXANADRoG
dc0BkgCLqh9Qe6EWayEZmCwDI6kmI4up5KaCsFOqNR1rQhg4DnxdvqnLbI1MGYt2391FnRjOinoC
TccexEelfKcdOg9nmChpRzcpHvxJNllnAKtnQi3Km8JBpy1h2coiawQfI0oKr8O8mxI28eb5H1vE
OKot+1Iy0ASIywdQnWgJv8wilr8W4KUr4duhWLQuL3Kkh9IgY8NGjRR/D070Tu844SZi9dUz+VNN
+QBFefi2mjvUZwgWbory2f8tosqQKS63DPiI5ezhjSJfZAgPVcRfDye+tV/Ul8ENaXlzc/x+7TDj
oKY16wxWSCxpdKdmVYvoP/rCGyAFGu+XNv0/hgK0RGZg6ih2jjdPmi0ZzWFbhCDs45eh9cDnzGwc
KesTKDowt1QXk+U8FJk0ApowC6oHaGCosvdx/x2TC2pMd2smI/2FeMlIa69XfNpVZkK40rtnYLlU
bTT1QQpQ8vMLfXldF1NYAtJYvNt6CmhSOTqPDJXqNXGfs/9V9aj+z11F++H7CC9y0H2fCEqu+dRY
t9hzjboUZks57yh1f30Bl8HITKc3Lw3IL2okBVN4PDu0X3h9P/11Ft3zOTgE3ppoZitT7cZSe1+H
vFMV+9VJZiN9XQCKhnh/IAAhqmXrc3rqnlo+xfy3LdBjjcsoUjlA/a8xMrHs/WqZ+itlPiuCSQtQ
xPJ7DIcZqqBuIqgdN0YH8jfeEDnEx0tUeMOnH+iWLxKebJaeM5wuASqVKM9z0WhTJY1WqoZIs2cm
M5s+qLso86H8oxtKpJjvu2pVtIKGY3IvhDv5OmcxjpqLh/K+lctgbBrZJo+7UxyvWDuYuQHMdGje
919lwSEAMsaMyB5lLUmVdOcMr/WBX/KwoOjJgWmmAIyMqpX2Nr+RITHlXgGSQbi/bsAXzH7OUeq6
RNRmv3EeSAW2JJWCepX56Fba+s9PqyhbJKXtjHe/JeiqRIPV0mpjGWmlKa6pxLnzKyZV1Zy2s+im
pMDdFWbD6jUvKM/+MOhaAfI4BKAwrCoGL52nV+yBJbKH9ykdSdAyzQhfhyW7YuLhRFWXK6XusUlU
1PykA98VX3LBljjeWudvgNLPij9fLAUC5+vmuHeYk9xQbKThrp7tQKn92xyffLQTOITF1eiAcZpd
7l868R5/uo64xqU2c/BnDoAtmzOwFbCZvQvVnpA3/3bEwAr/jezlggWapqilZQ4fkMPPm6PIzjBN
TYxZxYFspu5Jlzr7p/i2Qi2IfSLDkYSeOPj8UPVjaiWqdDKr0E+lGItQDG9IY9cFG9CvT+fWjlvZ
uDJsnAkRyYahUZKgDOjSdg1hxMBpa53vPLJB6/vAPUrX9tEj7auGVMoQxZL9Qgxgerof/2FigIW+
cJJrUzA9A5Nfjx0xKy5qCanjyTTSYKmzAVEAgyawIEPbfiLOWTNUvdwKWYHWkC1fb+QCiYMF/8bf
vV0xYSu+up+2AyStOsKm3zt7Myw37RSiruQhpGd1BAGuPNTjxLVVFf7lpHr1mRRmZpDNu/ZgaePE
BtZ68upYAWkygxUn/+OZMLSttNaMuiuxAKAdf6qcmtsMb2rZ2xM3HA9e5Dprr7elho70Z0PF/Dza
AdwsyJMrsuumForZX8DOWOAxPd7sUKc12z/naFj2BBgeJgQxohCBuzUfnFYQhpLxc0GQ8JdQjHrz
J5S2NGKPYdyjpfhc9H31ThzPA6CRaecNKYgCvVD/hziFRuAH/9G2OzZoTUPD6grxJUxz2csLO1LP
Eat+kpYStbvPuQWYzsuckYg7q25dVYkMo+v5YH2GzeuQBJn+t3Jtdt8nfcHSMxhi/DBv+9YoM4tW
i5M4H/ETNfZ3dAn5y8T4HDT0hsrYGQ+406YK3rfCzkwsAjAM3DlDJ0ivzHkeXbXhT/wwO4RUtR5d
Ta6AJ3FZqy5YatqnlSpFP8ERhbQk7yN2RTCyW77+M6Lz+mN03pWJxWJ0cUbaoMkfC4zjnwkNtQQ2
dL3aBKEl4Va9Fv4lcmH6n0g/o3y+bvnsQ/s0x+LyzzblprQdUmudDLl2ddZ6U4BTzLLnjHrZ6BhB
XA+AJG0Zs76Khde1mnZf9uIm0ZA/1WZZ3O331OsYF4RKfdCOUDYWzWFjO7c/XAIP/aJhbf8aFsYE
xLuc/AGkb85in+dboUXHOAYC5baog6P4KcmmyMzV/ZsqwjPVLkd2veYxfMljdiUWcBC7kRceyhno
2YF84Gm1xSgiPLXlTRVdts7DOSGjC9omN29Wx9GiiysG6kN7QoqfxFfYTBU865BFj40X8q9BJ1u0
K9bpwusTxbtOSHCcH0+MUOCpg+GPnXEs4x6NqIJ3KbaPuPeUzzpvH1bpRA2oAl7y9n1A/hSKOl7y
p/1lNLnYGjPAng35hNaX9SuxMrq53J+qfzek2jtPuPxlJvQJCeL8hu59UprFOtJWh7l10r+ZfIiO
0LltC4O0ZCHH+IpyAoMaDQ0NsBANsgVFol+146mMaxquoulYujEkrX0pNtJD9OeaQiH2A9zTfAPA
0RddytdVGOO0TdU3YkgRwxqVhBL88PxhNmtkl1BnCnaOQ4l/3mqVJl1ngbIIY8cjyNm1RjXPUXsK
WKM/QsEcJpyrQHScls+GGCEfxeXJbQH5dhvLa9rZCc1tYilgynSAO6MOSjMGXsnvNbHiGVYpjMkY
vsn5KeYIONgdzmgTeqp0xtemr5hiuf2Sfd88MU6taWivCmeYRIBcTeSs7hcgW7ZhF8ORJOvlbs3Q
TupnawJFtt3f4rqxJxfgJIyd7GUh3l99+Kwj5E7v9LLsD1jR1stbqUgvWHG4VOccoWVXLFs12G4C
EJHFj/pRalxJ7oH3L5rx801V+cpxMvvIyP9x3UWlzRGcc3Dj9ow43IMOYaqIzXJJoTksC94dT9cG
8auKdnnAXr17tjOSsc+INOCyoEZ5CbzvQ37mubXBE1/GiRUvZ3KoaML1sJA3jL/naLDHnPEyTycG
q+8JEMfJ3LE8AAIFg34dUhCpqU653J9iEMtmkg+WW4V4s2NUm7XzFJQgYXH1GqHd0QjmjYvLC1Mp
mGt5bI9N3/f+jp6M511EIyXw8yvRJ9WGt/05lMRexwQM0RbwBbt2h5D58FgO6jSkqsqbDw/wlMvf
BmEckeRPRueeUjUJyo5oxIYQDQUUAw80pbhrZ6pAAyxVmhZG4hHHbd0Cv80nyqD2uKcBrVLiRflx
XyFzoSWGkh9TZs0CJMGpsQHVxYCavriEwrtLeSa3yLx9yWCmPfcgouVWIRq9cfqU5LiZ4HB9ojia
zg80/ErN+Vl1hqyArdjz6GkR4DUP7xJ1WwKn46YFyMtZFcE+eEPw3hnfaScOI411WIlykeElBAqQ
8weyJd19MljNDw6028EGExz0rGaUKrY44OwnFln2o6K829/tzBZasmPWy2BTeUus6/Z8mMwI3y4x
9joZbc8UXCiVzLNMxJQ4p7ofQ2zhaZyycooIrb966l9OAZnCqaH9ID6bdcLneVZyJjWpXXHq3MAc
cqPyZnfSPgP2sJ1f98eAmqB+1lwngTe/mY4JBPIXaD3LrBXpKnZChdTr59sBHfoUt5l2nDO2QIt5
RMbkuU6E4NHJ4jAUtpu2OdTg0ypbQCm5FHfM+6yZ+I5CS+kN+Y19Z3VNNEYmXNxrNaatomf3PRbF
EICpq+14xrY3w1eTDSzg9ZjPbbzeb9uVxJGi4URPvsogfiof7fdaPL/1Sq1cNgT29ACJtj0JxBoC
jJtIJduUwKOrI9zBCmrNGxKgJIHeoJkKQTnaqWynxY+5Q11v9iq32yPeDfJdABopzlWmgMgdG3vc
YvKpgTmH/GnxxC4iJ/TU0DJeEG2HWM4dkNCUEBSIu6mENl9RKdr4zdZBgNXzDzOVVT1vG+sn3DVk
0W2XAzT64ZUzyx3Kr3i6DBlhEJ/DH3gXtgfzp4CPMi9ogfVqSk1XJjN6tGP6nHsD6EGPJo1tmUYy
6XizTQPNOgxZ0crL2fOKyW/2YVKwp5iRTHT0RE876tFiIfltFazbTLeMqWQBik9J3NSilwm2bZ4f
jui2eEARXj3G11dRDfKva//KTKjMsf+5OZXlFfQl6/49PlNiimxZvKmI46gxxKWNwqrD5BRZHPF4
L4m+Oezf0h43rVYGQDIKp0PTBuYGS0qzWa66kOEFeJCyNtWg+qSJc4KmTQ0Qlmh9fg7mAdzS6x7k
yX+WDQJpsL9XUXWFH8v7iIhBoWpY0qMRz9r0FLXrcvFCo0y00v/FhSFNmQISB+mh3TQdFRgiSyJa
kcgLdyUxDmu839h+VvKsZLFo6v4j8z8AyOshHJ9Id6VHY4zhfzHuiqqNkzo0tbBnOc6BTKNpwZvJ
umEdg0NEzuLzMfIg2/UOt+fYa5iZyNDa6TncE45AOKbfvhgXD4UNp6rvXFr46Wap0s36+TdGruv7
OhqELfU1rxTZWfg6tdW0Fd5E3oN58h0RJPuh9Q4LdBrlMd0c/OWbGrC59uZW9G6sBoQ3+H30cFEW
Smm7kqBSk6G9w8rVAtMAFGt04ptK+6uqBLCKADJlvpCgP9T/8ntJS2oB+Bw0F2kqeJARd4R2cElI
utCi0DeqcDz7qecb9n38C+Aycg/TKafhR6uQTdZGoyWFZfmS3arrwJkir9+7A97rWqNERqgnP92z
viT6VKAyiRuxjH6WwlNCrBK2f8gEl/H6q2/AnLbcRrSsPGKAJRZ1Yat4wc8oOygmsi+JTHuMJUqq
8g68j303D9vJqPhGt+diUgXk6RThTeOpqIQQEuHoiNxwmuPB1lT/HWo4hi5od9Rlsfe5WROl12RK
n8VupZo1CPMB36Kc24TGWsm7Zm9IiX15H51DgmjAMNYfRUrTlHM2gWOD7d/DkromxB6H5OPgzAj5
OwT1SBQ7gDQY+sF/eIlmhbV0+CrohCALffkBVdCvU5IFDqU4nw6YoNh5X8QX8JfiJp9+eItFORnH
c/CMhgJN4+jzV4by359mFELbf/1fPjCkXijgLrf9PtQBZPwFHL8AmSdbgRbo+6+yp6M0iBNxYN8t
3jgh6qcW9Y2NXfePacIsIsifQHkl9tjXW2PrRxdt1voNWr+vH88pN8NeuBu42Wz3lsU4xhf0+NJg
TrBvNOa2yiQSuKnZik/UMxKO3D+aLKaP/NbwXySlt5iT8XsBXt6YZeLa4FsWGkqQo3b+NMkToWDC
RqOS+8sNt2Pn1VQy5va0dDEP0LuNtqgDv3NP4h/PheOjhKVcXG8Pg11NcJuNJOQsGrQvaMgFBQpM
w7vVt0vEcbDPjeKAWYD0ENtGTfGWjstpz6+3/vBY78kurdhkA5wtou1+gErXvTwNf5tZLQtEa4yC
za1o+ss/KfyX3ogYZ8FFL0ydX5udg3VUCzf3CaDhOl9+XT0hV7TCRfRN3iddlAEqNsuXBY62Uyzd
pTXAnzMqMm5pK6mGFgxQ4So2qG3hHrmTiPZhBiYn/SiDBVHWP/Sy0xwj61x3EyXA7Yj+BZ5dnxYn
KCKNiGvEJlcRRdpP8OVPpWvMdcqI3qDdVBgGIuKqAMbPY617JZeIGXzLdo1KWvAyeHaZYqZFHD+K
gbeRGZE1E+Eed52okxsVgODYR8QhIQi1veFcoiUUKuI0aP8rcGgqRhFw8s6DPkzF0G6eFFCTzzGK
SZfLvFUfJgo669xy751XXkSU/tXUq8l2lbTMg3vp2yteHBZ2H73mvI/EmxF7lDId68j8O4zTpfvn
mNkhOD1/QNZNCh1/CGCmqSbvmUs7LQC61y7kTMunc5+dlxmVLGxvDkRRhLMFOY9qZPrU9wUqtgB5
GN+dGkC067xtIk6trj+FR6j0VlVIqGU+mo5KIoTeMNl9mBBbIU45pR4C/Fvi67Yp3QO3mG1ITP+A
ilPFLc3YbxkfP3WV+u2nZjq0lhhu1yK1vv8rxhwcl89Y0OqQy0K6BkfaIpd2rSRT5r0ku8AoBWBx
nhCLU+zMtXhq8KbAe5Fj+8pfFiaGb2IAh1xFsDMgjuQqL8DRL962HKn2yAzXHWtVL/w021B3nhYw
9BOomrvuE+vgEdXzEt7Kd1c/hPboDpR95mpAP/5rOxMUSOEuqzSPHEKAfxLw4WndduKPlTgha1q7
TKa1XQ92blO+ULVSHL6SlHtZvz7rt0HE1dYsv34aTuFUCLs9rfLxg6FdWFZ7DFKvHGylgdpTTg0E
vjzntW7BpoE6bEB7XxVzLveLB3D1cGkhLghkXXm0keRL9ze2akUduIguepO7vmNaCzL10rJMDXI/
W9Bqr/43cGmuf7GsCK2je+RLbTo0b8KyQmRZd3qEYAN9jJOdFxdTry558ALKlS9aNDmakdjl5Bx6
SD4PalvByXy+uILpw6+os4nccOSNFzLoKNWQjADryA9RdEQgYgCdRZ6rO3NzbdXHnPscQE1/K4aY
TrYRY+3w9egf7r0QVt+o5XXlPUsc+n7P7bM8asnj9uQIqDDYe7iOe31gvlJ2eEadvGtvCwz4OayO
yF1uoOLkibOFhvf1S6HQouS0vE0nX2V3hTDhsYlHnoQYerpH8WGw32A6Y/RGmCq5JqQc8P6jAahZ
/zgUvbxPW31UGqM4PdMNdfipMIlYT6vzL1gNLwuBS4wtS9bZ1rlQc7Og2GwlmWb+ckCPf6AdTuK+
oX05wSx2fE8sTVrsYgbt3O7y6VuA+1vaXWfioRctdGg9HTsQ0fVuZ3LerhTqZ2vTQhQWomwPv+hL
v1cqOfkpzM7pMddpBt2hIGxijjzkZ++jFOL8BIuhxL/NvDySkASlxWHFMvAiSOzDJJs7Nc0ygc5/
Tl1Vrk6ItqGLOKA2r5kebRyVxglGDCWShSLnStP+CdToUf3LLcT2/ZFwM0uHXCCc+Exsx4Y8O+n4
sTDMiyiBJsse1k/35WCz8rc6hFNw9wyh5c5g/TXFFF8Nc7OYh7Ik9qNAvBaEylhBErB8pPGX6Z97
vdGBsVSjHXXD+Np0MpiO8N2j7s59Kj3VihD97dJ3y9v7TYD3ZSTnt07LlItgrt5qJoaHJvZvUozX
CWkW4Z8l3l7EENIsuphAnUn2NwWrimtsDE7o3vcnI3iQI3G7XDvrHNwlgco4c24ot/BqmI+I3gXm
2Oj/2l6MvDn35SS7C2XN2E0XyGVkqRDcxbXlM76uPgfer/td0aTutXQJcgD7E5HBs/jpl9+bLvwL
ThVRgv6O11VWmZZL65l6U30ndzZQfU9QaX3iKqJEp1hQ9/mE9W1QNDBFGB5zMXh8CR2cIws/1ZVp
XxEMoOYujyyenavV6Pn33lLpu3ODhzdXjgj8yQuo37YeYDMXwcce3E0xhwEtC9GeqzD0qdz6C3Jq
Zx44ytRFdOU/z4S313gIbqhykZJDJpZZMCgsreX9QEWi99EY7FTwwG9NXIQ9oN67RtV/WoYVl7Id
VNFHHN+EpMEuhenLXh/xp7+0ys93W/BiQgT86K5OTQLGlfPawUR8W8YJQktRsuhK7hT6bMJ1ZT53
vLpKUq9VjOXfdggwpwlAt1+ArV+EOHQghv2oZ5Wucg1JE4vVtRLjf+5UAEHj64mW8CilXerYLeVp
BHGSO8cqzaogu7i/Ed7W2MBbgIIpoT9DLvA3FvnXfHC/XGRwk8+004HCpk7HCcxL2kxxrMsJm6mY
JQJPsQVD7gUZiuQBsX68au5nX6UBSmR+mWmIFMj3wsAs9dneg0YnxCOdWljnbTiH9xq1Mroxe6gY
dPaHguduiHpyxx2SJoiAwYqHUKQUFzVWY/yhkhyRONP0L6y1OfBon2BRJlQjV1QVcUl4bZ3s6VlR
tpx48LIozc9o8ne/zq9/A5IN8EUB9KeuhEke7uSGSkRf/UqYSDHESNeHb4D6oKfM8DOvnKuiOC0c
xzmX3rn170GnDayomFR+GZITJ/irJI8F3rKaL7GrX2kDEuw+U/Dn/dxx+WCE882WbZ5Rp4JWEJxb
bxShcGXFsBg/H+sgFCLlvwxA/6qQyo9/yNdiXWo+7fJyzSeODwOEGeNDTIrz5RwAKdaFoyQdnun6
otn+EYOrgwhuPsThUkeZ87aVSomDdKtN3J1VtNKipGJdBDSPCF/2jzr4t45ImA+z6f2CAuxGadij
090IrWbItTBY32NGvvVU982Um7oA/4yLTHebkGpBu8yl0X/vSL3p91pFHRombjwaKawtLdbRdqB7
MVundVsQWlYHiCac+CSBlkIdFsoebaT734mTbt70g8pCYoGzCfLxIi9mPePUdnTqsq8XKRp/Y1o0
nGueMhD6qUBx4wML+FfyvzvKthsNgUX9QbF9o599N0m7Bi3W38TaJL252ryyWS8N9wXx2ADHtnIR
z7FYJcHJzfS7oxPWlAnLhEl5VWkKsxOQ/iosKluSTSF23kXcCYX69iYqlNuX6dBlQvuVy9V7O1XV
qvCZYx0sjHJ1nTkg0rLS1s1d0Fgxa/wS8SPL5AEH5GkYT1b24i8qwdC4vFQjkYROZO2uWUalTsHo
vxp0CEKS8jOBL6000EtgcT75OvagAsjSzy5tF8DIugRN3KnzRxgCtxdz9vuYBpmrrggFIz5psxJA
Qi9VQpXUBns1b9SiZwIJORgyLh5H1tylHYmlA7Id83OlovDxeBrCTVBUoAyxZdfp55dWtU3JGuZT
7xyiJ/MB9uCpY0zBLV5xkKngpzQYpZOE0Rlwd6TueZe2nKO5pYCxM+Sk8QfqDwKZEMS4Kn3Q7hqL
Ss5qm08Nsfon7DZbzsSVynWDT0or3JerQ0KL6TLhtPTDnf0XqscDerxztBcYOP5ibm3kFC60aqsh
51HsR5nlIVC13i72Op6rOS+uT9oPNBy3LqneoaitSX3Q4JlsRrmjnNPw4VCH44eeQCA/vuL6LilK
TYjWrWSaf9DwPTVZRXEhUezRiBX4BtNqpy8aIFEprljR5s0IjE1UYnOOpDmvLlpfRk0cO5H+3cfE
Jbnz77V+nJZcnXcBHG6mOfrbyRBJwFFsjc+aIsV47SUgGHKTThzt2uk9UT0mJ0BfQiMcWDy0Xinw
qf7L1BULyBV53i0cfJk9b9ZcVfejUwt3IpuKNSeWUOKtFYqT6qtXsyNPiAir0IHy4rcWqwVnfX1p
yOf4U0TRe1AklfsCY87Tl9TjJDEJdIzD4WWvHHGuqMC2+tRvIg3YnNkiK8XtjfFxh13NmCrxtsPJ
wYMwZX37UvO/Wx4hcEUeYzVLYAteboqKxCXqVTqrnXhI+Gcu3ZcTPlqYcoo4jsFW+mOKEfm/aD+z
IXRWMfRH1CrqzrHeju6P18lCtYZfFTpPLFfQTZXkPGHiOnGhHpRln7QZqpoYJR41lok6Ftxq35NG
ezIXWm4Sk49quIuqDeeNHS5BsGoq+EMhBudvvf6L1ozcKFd4plrg9SxSnXVu1IXCPYG4nMET9fDS
nsKl031DdXIBWpO06WId/8ypqMYC0i4aF/Ff8oi9i3QVGuDyA9KdIBCcbhMXUa9YS5A1rI8OI+rI
cPC8hGVkgPK53IynBVu4kF+JraeBPfbpUSDfyrctVrPRGQMXZcNUZUXWVJHWxuWkBLN/ZK1RWqjg
OvreeyPKArfjUAdDuzRrydWkryQsNy7vqnjXX4262Af54v1f356EqME9HIcoLlJjdmn4Y+NPoC/8
W3NClBfl79e7hhAt26+HnKOYeKzz/+i25v4/qynaQ5SF+0VvWq5/BI6IHOlDqIOzUfZm0x3x0nth
UnBVzTHcvoIN6n4BarZpiLoUvuZOO1c/UMoOT5zeljQ+5kdT9/etOVlwruqJ22FjFPY4Rhur4Yw2
a6KgYhHTRA5qhpIkRYNeEZXOtMhF7/0J0IYwD2yjkOAFYTV6X6g9lrhtGIh2nYnWEDzZmKiNV6YV
H/xhJX3KP1j0JwP07yqPJl7MsaZ7Fr+Ddk9+Kj90rQ2rZvNTG/HB4JYNzNBE4/1oCPkSVdnQcU5g
fqQrrnTAOkmsHPXWy+ZThmU+pc+ZFYl4Z9TRdhlYNDhSzboAvQ07aFh/ZUSomSj8155VWT4s/8CN
sTla1K3gdJU+o9UxVmayWJJInTwZ2kp8pVxC1knbxH7/qTobd8dKoG6/d6mWl/6WJIipUdz+A6jp
EqPXxk8iLvlCwr9Y5IVMcyCnyLIwzPv+x3p98Z4OugEsVOjvSoEKO3/My2KBpyxYHvo3tEHp1r++
pxrfqgWM8G3OfPEY1npZUsXgGw2YKedc33xz4XPAbQIxn39KBEDZY8r6O7EuWOxq77go6NufWsbb
trmr+QW4DehV2s7xv7V7++69EvDUBsjLz2d0lJViudA+85y/LkicjJk0847NGMol8DBa82zB4JT+
A1NESekTyPQ0ydCLZV1HSbCuO+MlzEVYvUHKoB9yPV0CDk5TKEX/idKowfqq+7HSYACstQHkOCrc
sntWvDoqtbGoYBkUNx2o2xEVI8DdMOI7ue676h0q8SDqgvGvvluT3oOjpftlEwBLr/c3bDhrmevR
rOOfRPJpNxZI4ICyrQ1ecREgL/11fqJhLvmv/DGEKOYw3VClv/t4fWNak4GJDi1LJbBWQP3OAor8
mW3LG+KDSRfKpB6QF5hQQRU37/0qTrTMit2214VQ9yHQmLMC1UynACt8zA5tWO83voymUF0kPJMn
uOxSDQLVE+ge5GLVnO+sIq/pzIP86gk/Rc0apIqfMereawkqZoUj1Qe9IsU2jH5jPCIS9MMs3tPn
Vou/IYjOT+38SCnh8uUfRIkNnYNZoTgohLOFNFWepdDiz4bzTzZ1Vl43AORbdr1+X0k0M8TedZaQ
RtH/wCy5YKFHe2vSgB0m+pChapGk0iwcfNlxWcyq+ZEK/ejXFKYElVs2uo6U8rvrb7VqQycD8ID+
5/PZXBVMWHjNEtGNTfqDzz2BYlzOcdt2E4JEjewJx1pD3UnJyuYg31FZ8kOObXV82XJGz2ysNmIS
Qa8XcfrkXYuB+A6uApnSCMFWWYloP1tJlVkySc1AIQqHYP/bTVr/tu70MPAFs6RzGSRjCqFPnSgM
IVKhl4g9VODipi/fIvTS9KJHMUJ0WA5o8Sgm/TOJqyqiadTvSq7TprCjYxEzqHVaaTd/ceJJu0Nj
W/z6BiI6vyVqbw4arLt0P1Qay7mwCwm7VJu5kyZeSJJn2BLxDac5pqjq6FzJ5MUULt/MdJyGRooE
nu71Fn08jJT57EFOqGs7/UPbdoMrAKAnDQGc4BTXKcX+Tpb3FirjnqHZKMOVgJ1ON8jifDN+Ted/
7/AGpuqyZOzo6qgBXYd5EizfQX5v+qLZegxd2tEU+78zbE6nrdHoGfC6sZuU5WauYKwcfh0lvmgC
i/5eYqD4R0B6qVCrsjU8ECrkhiY80dM3P/G9RXrovcnZoD0zwGUuPuR5/m374UidBlLOjwwDKDy/
4E/OCEDln+tH3H16es/CWJDkK4wPXlO/VoukFGyseM0DQucIZM94F1fdgD2J9EI5W2eyXAjmsCdh
qJdz4HCexPKBcyE/IEs8F2QppFrudT19jW0JxhUlqa4CAny8eILxFQQlyaXMB2hdTZWpywQhHRyv
X9uXM7IfAtSoaWbJQKfTj++QdSjpzgZhvH9ihg0aR/NW0O3SLik8xn76dmAhSpEDJQt3+3k1eJ6v
/hNXguQIr+suQLt3Our4NhJcImXCR2nvWG7UxaKJXulSFyPkE29GAReDL7uxlQ2JjyA6gCqwr8Zw
KQUg1iPXFVIRywmNvOKLrhrcTVNpc67fzIbtjZUaNdeFtBPTWtbouAx0YfVxusZuUaP9qFHCH5q2
wFQo2jM9yBMx8a+RI/clPlFQDmsnVb3E9H9JNL/vEh6rLG3KrNYqwN+fHC0/TnH+o3QcB7cwQJ6T
WnOkI91NVRolYGLt72glhde6f72r7moKG7OWhzeU4wjr8QvOwnF0PQwn1eB/DCSqoycF+oA/jocR
Scgsb/oCUg2EpPEn4WG+nXednXR7jhArWUDJBy6Oeult5sQZxXQkz6tF8zNs7xXtl+bN7L1iSHmF
BWBMoicY4czH2Dwi4xyO0Cl/1/6UtlLvVQ+YsRHfA2CjEwTALCxowqlq4DxukbC10p3wm3SYGoAT
9Yv4bfe/tRPBgMievPSsQ/fvryAA2Zq7JReNzQugdCSDU0yDR4Y1BvsmujcZC9KUrrh7r88cnvPi
rdXCnJ0WeO8Ciqia+M3kODhavYMsZVP+S8qmH/ivniZYrixXb3ag/9txwbEaTQdWYamWflJ9PIt3
j0xI7/waBV1grZk8xYIAHTp92bgsKIFxzjCpI6gZWCnb/tfT4dIQJzZC24lawoS/oHQQUsTPk96R
RPeAAPV6o/xBhw7zeV1G1v0HPGPqcR7BYUuKOz5fJO4ufi2uBKClk001Y0auS4rpUj2R2OSDXaH+
zd8l4rzOuLiUsIBHbC21qS9ekJ/mG1tLpirh/HDoYFgNF4eMsQ0vrX1ABeCK9cnpKt2F3w+lmX+7
6zuRv3cPsjrL+oK2dpRCtwm8/PqMZEQqPEZCifsjV49VI9yO9O0rlqx5ZCzEjF5zw75RA/TrkprL
j8QyTdi+z+gL7NvBOtb52FaEGe/eGi9nAgg2Zea+G1jLep1Mlat5cUdc7RxTefCiWb1wnnlBnD9m
TkNJ42jwoxAJkrcNiUaCN3hN4/sY8+3TSp5PK81hrP/9khWm9sgRVKAuNGvHT+ly3VsE4co/iPLv
iFLPXBFn9EszqpKq9TFsQu2I+I3ydS3VBHKslcM7uEbc40JzdDlkp24ZLrvSz+kxADbRT3CY/4UZ
bhXv6k0zbtE0u21wfCe0MfGrBFSPevkih5c57O75EJal0wdfJv6I1eR7/eI8vSZwU2cTIokm0bKN
7D9BT0lxJu6u5uxq58kPfA7n/Ro7J3B+4XqSbiyH8shX6vCWVJlqUPujxC1DjblGulASyqshvoo2
8/O/M7Yke6RJEHsq0yUEVCoKiBaBMO3LdxweaAqKb3EU1LG/pL2UqRjJovVPhPfQEhJagZp7aQST
4B5b9QWjN0hM6wwDXVMuk9Vq/BVZFWKSyhFGuGfMVZWdGRicm0MCegRkdSZKSmIcsyog2IoVPIL7
iIUdjfw1Wuw1Gz2eh/QwUBb1ycJ8sGZ2A9vK5PDKblEyukXHy02YeK43unBzoJG+MLkwQFGRWFYS
PUBzhg3+uenczONgJiaogMeGmV9eORpNCHCdW0JFZ1xzyMyBb4G96oGunUeNzH2moWRtuDpJql6M
/X8SF/Wqf3VsxaFUzAj8TwW8s8TMZiN9lD64I+uw3Vi8OcPamYZvK9sTzHKomjrKZFYToNC6NXmy
8nSckVIhKHPsYNu7jLWP08mAWUqaBFjz70L2BkMojRuLm0rJ+gWSU5Ll1ozxBhlV9Nt8ROwOA20i
xb0Bwdw6rWcldwdYgMrmWnTiBkmTKivcMZw7i7Qr4KSSvsjkgR1ClDZbv/ZdJvYClQF5tyf89v/e
Q24+5YdoftYt7px3TFy7khhHqXpAF9/yYGwTUe2cxSR2q7oSmzDN+/IrUhXcf/DlIADHtKfudIsW
0xjuKistzyg0Zh1uAuzZGSOgafO/9HIp7AE0w9GUmU1w+vuEw0aM6h4zOVry8uXGDZfq8SHb1MSI
xc0LncB0zvSw8V2gdLKUV6HegWD3BvRiLHjvxSS4XTexM7KVLVZf9ShwRcchJvIk4WhASBgzM4Tj
tmC0RJqeQj8COR2KkWo1hgwcMPAYD89aiMwT3PgzZe126S9Ky9p79I8bY4obsGnG7Z03zduBPHXQ
xVDAYeV6RD1EosE90694pJM+zYy58U69rks5TxaSUFFV1voHU2mCOqjWoAnY7YZtFejtQGARQ3vy
wOeGKuf6BGXbUAKA5IWdNYyNgrRIP/nD+ofVoYQCdWLMJ0fz/gqaW0hcuGrPmxObrmSSnLqP0IAG
lCP7KCTme0eFIVia9BsoYNaSnTt0ioyqTVoUZ6RQ9MoVElmSPrILnmyFhPZ0GS0komagszvhsk7k
ioOU4gbfhfm09gXI5bZmLCLmbsXV6SF8WsB6kQLA9MIpZml9VQKVeMxMoZRqWjAKGWr3uuMmN2Zq
OgIc5K+fSDbAXJ6AQnZUKYMy2keGtsTclaHr4qLxN+Cfcz6fEF1JUiGwJr/Ja3sA3XtaP11Mn0h8
0dTB9VpYuWKjF/1Kil8bOcNZbMFIX59LqyVr8lqxWl8619VXSrNtWeNuA1TDzSSUbqLXReQ3nONH
pT/JtG2SiKswLWy7Uo1BDu0JKk8oWhY2qk9GSosSezwY1T51sXPoGTbHwZz0I8p5CJjxLztmzWbT
WQ5QRS3Svgw0Z6NV71ZD2x++jAyDSejyhinR7b+ZWGcl8ecj5seGrXQlv1+g11TotgfdG2Qm9/za
xdqk6ctdO9Vxc2Q4dgJXHVRUK353g6M44TD82y3wGynyJSzgR7KW1QyJylhAA8p1wHEyrmI/liWt
wz1vJhl6lHXlhsE49qZfesho+Xn9vGSCHYD6hLapJb/VJAhPImXvA5LCap4+aCpj71YMkHWTxK/h
r2zG2pOzaUwAlJ0ec9Chx6qpzXBGA3OUIPusoCC4PNiZOrI9Dp7jv7hNsNpFxbrRUvBfkv/9P/8l
4L50pzMQxYnqUQ5xNGCVf/R3IkxjSo8lYpK4hcjXQWu5LCcGZNB/SQOEvZsdpRPVIT0oZFXqLDHk
OtIyPoAY9waaAdWPhSzIsm4VWolfCWogxwdXzFulR2iVjTfqMW7h8QEIVbuZCbEW55AAuXHXeP6Q
ixKneKPj83XwiF7iDtq01ZA4MPfBqzhv+Bhmjkr8LOp+Bc5j7NARMOl0JxvdzTW5LGP3kZv2e07k
FPT/oOOi5kkZ3AFJd+IWfF6/pLz7BVRafkDL0K+IopPW+Yii8MS0wOKcOFcO2eneVMWSqcB85kle
8fXk5TEGAaS6ibA3yeS7T6iKSZhEHGgqFTUQBGvV+lhR591E8Or6FjNRuso0Wzyb+7AJ/JEbCJd5
dSIQKFCWvdyVsPIy97udRVkiUOmWEHNp8op1NzoBaMOa5SFUrn0Oaai/qFFziiCprilxuKMcU5Xj
fnpNBMJ/K921YR7FwueyJBZAr8z3e9ilnc+34T7HZI7Rj8kOVPoc2VClHX6TYFBXVx7kAz3LNU2H
aO9+19DHv0s92T6QMCtewNiwMRwSSuUL3dQzwzdseMbINMVpOy2wvctAHl759u5Wu1fYWbyy12fO
8hvYThM+XESL86gW+EuKeSUuhQEDH5H6eEdmoyQV113OvJT/RtS6G6NDiGNMi1ie0JzVzO7wiig+
eHZjKXN57pl4h4gR1epRx0AgjQtwVEM8pcOegFZn7dFJRv4kpML1uYYBmqcPmz3b4nG/5TeftLpA
Wut8vIfhaja1JaxVG3QTx/tz4nzY6oIZ/trW+3fccsWNqKvd5Df0u07SqmgLUSHjmT+jj4wTMkZ9
NRn81qM1D3+5YAM8WfBMlk6nfz5MmGELHeMRceMBAW3G425070O0173jQmWbCkVWXadsGbvawLgI
KhVGKVAcjXbSeyMSsLRdN+AUvKToZFIeWuyDtc+dItdHUP2SvXR/+P6z28DZthbyWXkIueloRtK0
LfNsLZcE0g/5e6wzRYBtW02RSXF41l1Tnrku90vhf8rgskfJiI8hy+9GZjtZpxlgczjGtsMdmYRh
QM1xkm/qHTU3MExOwQSjs/ApvJb5A/QJedOJT1WlcPygdcbcr0mK9dgCllixkiKD6BaYa5osw+QF
iRMF9oJo6qCvPWc17OiVVOZ5b2F+b4INLuYAW5kePRqAeSpeDbHSlA+UnICbOL7m5QpCk94otD/B
7bz2SVYTPPApH/xLfQFdlE//aycfNvojXDGw6Ew2ipPrK6WUdXD7kgrmRa0FX9coLm5OoZSJFVCe
geBYHOzm4R24PBnPcbKyxsZdOTwY1HkIuSH1E7sry4+Dwq9zvpdGVAALkdPqatD0MIsscac1p0va
qPT8CkVRrU/FYkX23RScofte+tKpR/LOIsd0Uk9U4V7bV5NS81IpKMIMOG273xqgEzQ8X+wkMDTY
tRJwJgH78UbEpfeMhAl7YwNLbAV27DVTAbPu7NKOZnbqNy9sYjf6x1dBWKHbZDqf2AULxPAGrdoh
zS8Z7f7AxXJXslokY0xdbDUOPpv6IEDNGtUnNtOXc0wH+6kT6IxsO9naUk+ED4N0gdtt7S6GDZNq
YDAfH7whyPwIwbfkac8Ch9v+dEBBIH9PS5Ic6X5+zeRZumjAtJ5C38cPr9xJKiF5KpyNOFnZA6Ri
pZAMlEfuK0yOGU3t1CZa3jc4ISTZEXfhF27eeu4BEbcwaGYyr6/2d99Z/0lOqOBrABRshxc25dpq
D+36Sjspie4NtY2e5/axK9+KCTApMpW20CqKDPBVE/5UQjH6sFE6u8U3thueiF1q3MJmPEAnFwCY
8nZlQYPP2gjYQozlF7wh/xdDOJ9MpOXMs1+7RStSSGrjsyrRUweDQ89Y8vdczNPLUt7bL74kTSNf
ehr8OaQFKhxnAtAusDuzFrT+UixuMro08/TnXeHwGxbnsmtM+dTrRbZ1dAD77LV9+mpg3qQNjXOJ
lgVzM2JtAYVY+cGos0D+7ieSmbomY/WPkF40VZWNZz4dFlVhVSI1DZABRf4gRxuPm8X1B6gAcQA+
YruzLT2Pje1jJndpiOiGGy4SUvH/JZCUJGj0IS0JtZDjdVkyfS4HNIQFwH1AWVA7ChjcXGc0Rfvy
hfxP/NjAInmMPW2u3wjsXjEG1vuPMCzN/O0axwpODnC6Gzppdd5aLjIb5rMm5ENqO2Qe8p3wcE4U
xWY45AicLB+NSEvktCvH4DZDh8fN3v5pyt22j8DddUoPy1HBAxcvaIdbwy4iWgoTzQmFWgGdOuzO
ZnAXbCMN+7bvQiETzWo/ua0GPp5hCFOiHuUjp38w1JuDw7O4Y/pXKwIXPIQYeaI6+BfNmiUEqbhf
WY4NkZsrBvqNLa6rj5LU78pZ+v/HtnZhjhGSF0uHwmbQvsSM0a9QNXQtdynnpvAWn834gLX3kazV
m4bxU/ufqZcSIrkrvxtAGxfEN24mz8aDo/tlmXCpJEX9vsKuZcO/vcnXk1pWpdtc6NbyuqyDY6eg
qka1fxPoXSRH36A1WkF5HHMGwKvb0d+HvSwEjlC0VPTGhhAUEPICKZVwACACVqrGYC/GRZolf2qa
3FZUCT/otAOayY0tDrqsXONd+mHR5mLoBpFLQGB4bfMt2QiMHmgPZKZOVhWMpzrURxl2dY0wOMZU
j0p5CUYDyX8gF+1p3LxJ5qkiWHwVzVrSTNZgRnY3ua13KWiKMs4zgBnlYfpdVmoYWeIMessg6S6u
WFiKpvks18GXbPj2Pjkp+pEC01AaYx+X8zIP9GMPo0i0Id71vZDFnrNIsSHIeKrDdHNR0nqrP8he
zzBTLHE0wj53952ElYKxDL6mEiAnHYbeWBZtDcfw1SemF202CBY/HFsisBMK5JnnkwMScSWCA9kA
7hCS2qoE8MFUPvGZ0nHrAIUSW/Fv4Y5SjNMLAFxYROJkQYvuKapIRkCX99HPHkAIpsCvXVvs55yT
2Ew18o5Ii1AfMxEBYa0Hazqg9jUlp5iaAHR7P1vQS2bXtIShUVIWcmaPTR7YLmejp+2J25FEMRWm
mMOdLTVd51NUbvdNYB0/fPBeRiz/uA0tx2jivUYhLZf1y75ZleiTh1NcldEqmqlzn5xO02wqxIc+
OoDelBFiyrGfy2YZa+D+KE8G0nOaPYVsg7aTqu7x7j/KnSUdT/6yR1swX1tdtRltspE5MtmW/6aJ
f3hzUUn1EvbPmxTFaIQTzPnSYrFnHZq2Scx/BCwkdgdtlB5wrlrLkbp249BVXUlr+728ILxlhsWP
2xhZI/boJFuTVHmnn+x9odDnIShcNYyIvWj1ZFhYL27cLak8pg4G5HZGuHd4gCjy5liESQuU0PQi
efqEMXDb8+S4nc2PyljzyuMmzFcieQfADJSopgEaG7qr0hr3gIefrLGWIxaoHkwHHL2WaBZ3XAGE
H0QO7Dbm9XCN36DMIjnOZh5gptacObqHsP8VSveEwpHw4J2dJvMzNDpYA1Vy/SfnU0Y5jWeNafzf
6v4+fxsBovHIagXDV07In18pK1DKBZloP3e6493yWbxoeNi8Qe19hUBYAfx9TPtiqIvMQV93M4i9
dxP4iFUHXU3ElvAPagemfbl5ODW0I+d/bMqg9JQSTrVKhv6hdjgme+KnOy5k/Ign7PFXEhmbp/T3
J6wH5yY5rfJllHUvdM2HbbNrJIr53d5uIxNIWxdZFoh7OJ7kv0NI0mzULYRHL0gdLqucxWQfAJuh
dCfqdeHLvLbUN9uku3FSuYd38WVE/Os4oJ3bNip/9Gytj0OSBkWpWuJFkEHWDwM/FBgK4Kwdqd9H
UbEoW10DJGlZhsoapxbD9G2nJ1Lru9AKQM7V14S5guDqik+eGdTLTDUJnTqFOyBRH24+BH2/0HQv
QY6ppGtU/Wwq16jq8X0zZzxigZrlPk0Y5QsqZZ+RBEuupWuAzvA6LU1XrztiPi9z/rY1izyH1gKO
+uVtbSlW2Hjb1D04BUxyoTJ9bJp1KsD3Qlln+myy8tXEBRPepjaJfuwcOMxl1cqT2aNgRwy6/4bH
FwAiDgIdjpN4lOBPraoDtNVH9J8jhk+XXtqVg+ZeQLldnLP6buMCWO00Scjo1QT3P0A7Vb6fVt4F
+yB6HtC9+kw85WJJkOA7MXHSslt01AhFrPU4y7We1ouwefGTq7MPkFlSLmypWDydrXtfNNzpOvl7
NURL1yU806UlprNld2OhsUOFnMr/WxhYN86yZ3ZFHMzAYOBvCw5VmQiO4aOjyUcvQ9gJTyezd99y
tvuqweI9ib4qwmNppW95m+qQYQTVRwp7XfNXQEj886zrTTklp7XOUfaFUEy6DPM4Zaz5AWxx0kbW
5mBjAGjy3JIrBAwH+XZ/nE7g4h+YzQ3M14NYtl9V7q7JHWrJ5D6TX/BxmtiryT4WtE97o8tKIIe8
LK6sVpTX8a1SYEpDxpHtjxRLQnrCSVS2wEtbtxWMHirMaKe5P69ioChe4rZaxzA04dB8zMpbeAse
W0UHtGj/tR2iH0mA+PAtIbZK5gxEQeZJnT4VPLWK/ILw8WaUgtWTdDi1CXDKbcieYCixgibHIBrP
jcNk91VNByXrz8tCuJaivMHSvEDo1+d4xl35f2si8Hf6pTv1voCl4NIwKbGYds7qa3rQkF0+1Q5D
LzoBKmgHjUhs37a/P8UjLBCpNancDNSjKu/zvFTuRs4jRdv+7QIf2GnCgiamPJOrz9wmonaOpjSY
9oo2essZ1UOR6qXHmdWG5xoqetycbI65eiTSRyRkScy4Vf61kjUux/eV84FjFUDQ44xwWLQb7D0U
Go406sfVIK9u4721uIbdh1DpJP0hgov760HRgGIGIPpq41NKHO3pbYptcetpTz8/dXCNCthMOxfZ
MRLA+y7HTkw6bUmBVGMAoxyVC+YPYoQpFtF119aTHucHaXLBSp8z+RA8iqLeDvPKtcKz9ldm2fvn
tC/88m00k4E/Wuv/zoCpchGANAVR5sJaedHWit7zXqcBigM3zlRdt/Vdel6Ha5NQPgnkNOhIiMle
OvotTXgwNR3dYHkITPV8Adg9IDrqBtSKhd8hFGggZff1kdmrSuSC9BypxYSRDXdHlhEhzltvjoIh
G9HMWDgm4tqd2laMW5T43U9mIwtti+4tvmAqCFrL28iMQbGnmYK7pLr/mHqDYnecNTdcNJ5TZ793
y3BjBzCcm29NsOZaUACVUGpqC66GO3vzV+GaRACs2Rk7ZMo/QVPwkYVJARrGF1YLUeQ3LmBBHdG1
C9mJCbH4eMDcjSB33k4yodVrGBh9BudIjA/xi51PoRiiRuy7xPpQXNirgUTlzi964dO/ktIbfURm
jQ+TnOHUUx4PsiYNfB2gpmiP00TmOgJXsDKcku8zChiODSLtRLU8BtScV73v86jP+o11sZqKjxfP
Yi1KbDNtOx8FPPwNH1p+7FakjBm4km6gQ0jGT07BcOz1qwoltEgs4qNnuTz21hgRRkv174amJ6i5
BduCU/5XD7j4lgi+9XVRvdMFhP1iQgyGu3P2d0FCHbUA1gg3qDeRxezMspXmwztiyorThfdECWax
l95WaWLq/Z7nBGZV+eetYnK0vWXBPmKvm/iE/vMWUtwRdSilEGXeuDeBwHcFaY4kGkGVYc0gNpV5
lj//8xmFaLPosJsp4Icis0W1ggTBbX7AWpwJ9a2uvcZ6hOVeSJdcAH967zE4OQfTE5hCQL0gXti6
LuNj9VYSTFlMO3OFg80efhAvlyyd3U9VLvu8TK9JSj0KF997OjXVLC6sP4sVASyUX1IZ6W8+1fpv
mwPhZXFtq0p/H06ks362VF0pUIco3C9kJ7FoxlhGlbu6Q2TAiRw2xNgn+B4cwiKLV+mgPthQ4Ghj
8tw1B4qlBpR3Eymcr+8p0HWZ5+8mWxEBDmLGGQL0sJVP03Xt2MJBVYweJ6/fYqirp30l/fLhoW5w
c4KfX2DyCAB82WAVLbFJb8FLFpFzq2/iNJHM9YVqRiZ0M/X305Al3q7PTRntdqj631RMla40eIUx
uhTxjZoezY/miW0z7I9/olI6PmQGzPaztW0xkvfKmNP2+zXeaXG4wahdWF4IMbiG42GtAep8ecsD
RY5hh8u/kzDjYej1JrP0NFeXTHK/bM+b5bwAl45miNBpXA3AqFRt9AW/I1+yvAok26+3GCFvPpZ7
dX51iLp8LwR1z9vQkBv+92XabJ5NdN2mDEX2rb5tTapkjgQqSO2Jq91hgEepPw8d8z3Ancc2WmMi
bbtDAIxWRRyaLw/oZSmLrQ1GRmKeZjLcux65tqmc/zQWoLgYSE3i2MdGvec3KLKsMCu57cP5Fl0s
pKIxSdp585fXeiTUsc//RCDzFA6uPhowMQABAjZikdYLawb/WIXAL3Lp8UYVXMz+cNx7U6nNLu3J
kVEqJMhQQW2LVjUQulKc4NcuzuYEArzcA5JoZ5TsHzgJapENpnYBQSESYM7BibZXpNBnJvFWR0iv
gJBrAbsQ93rJVKgK1m9Y1fEQ1BygxixXnj8VRtKtAOwxDZDKDx5vFTj0m81wIOKdFGwXzvFAQlfl
RDpCYxPqZCiH6IlEQn9R9Hq1RAO/xQbXGweT3/Kqd0qfX6y7mLj+WwS0bIJW+kylaiStNd9rHSTf
uvE5rmDwfLrg2ZtDokeaEJp2IjvMU4J4LrpTt572KUee+3zTnTBjGu/DYOmLubODdhXjxkLNrAfQ
xXh0gqKzqvY2+pTp3MXTWJV+QTVcNLv1YXWlJ/zZ6ymYGo9jGqfTBVzqSMtvKDVucJ1esfAeaHRn
0Jx0kbo6DMWaGGFYlzHO7HBZX60apEuSyglL7ZJkWxTb0vI1QgRBf4zzylixi+ThR4jFK0ss90Fo
u41WqZk5ZnwyJei5OhHH1/ItA+X8iG3HGKVQ7Qi6nkW0hfhSx5iuPvnDlmZGGqG4pcHc4l+XPxxK
yWTSK34+Giv/dv+X59EtTZ8HcWIIYbX3FPYF3U+/t7mv1uYqFW6BB2padAj0NEZY5OM3DTy8t7uU
vV3v5FAiUfxS3UYcoZ4GI+ABgQoloOP0d/D4IByKacfRA0OVzao5lY1W5WbLJ28AiB9E77ghYPJ1
yiP3nFnWOY7nc23jYtINHYHxXxLtEd3Wzb0n6rpNj4mITkmhF9Z1pdxl43zJoghq23PWAYXFN876
MF5Uusy8roESpM+2ozBnNUJ/1H+Iut8l9fK/T39o1FQ5cOeaZIpNhmJfAbrl2fZzqoQ1vqrLtZIU
UfKLxKcfBPbP3PZboa28q/G64hdX4exvDLLRiLzCetM2IpKmWBEyXgts8FqkKNDCQSgjiAH+lPQb
MwdWY/VzhFunsWbWjjT1gNWzf9uX3AZzGF/1dYvy5MSr8cyNTjq7d4n0wwZJ9TeFGGnVhMt84BrM
EprWySFc1QJw17rlPx8j640LmvIszBTxykZz7/1awJReGazSwgJx+Ju7FsSbZhcpNSPCQzsG2uDw
rzJJyISLGgK7vPA/yB5cCkd1ZelgebwH3REe+b/b9ht9ULskitXUjPamF0iwmpVTlbmG6fUYPiUL
TpZVeOr86n5z8w/4EbozK+ri6MdkD7jjxLawMX+jIYeLPaT8Tvrm8b9qHMAMNvmAMsjbhukcg2gl
Z8sj44ebN+RvuWW5wjp1k4KRe4hlmQMsE15jAeYAlf9ug6Jx7FvynYcdpTKlCw0RMpvViVfCwhMJ
kAWAI4T7QY/XM46Lkok3nuLHahqUxlEc4mnI8DVQb3NHjTbo52OV/EwxpRr3/68qUHKpHcGk5D17
AYvLzaBJtpkOxuLUcZL+/Nu7LKCzJ0RY5mXB8AFxaIDZzUNDCktQKwV/vj/FBbOaR2T5qsmCPmjA
gKuleVOk6vfQ8F3ACcfherJSrgunIm53xRjJIVqUyaq0HGtFkfFpKMs5VmQnbnG1QV+Lf4v7waM6
BhnnbOphi4G/pPL89P5Y8nSdTEQ2DBQPdJ65lwdYyIi4EKadg+P/FBjf0tgPk/zkLoPmAoWp29Rl
9Hrzqwb2tDg+EQwV+kP2eyqfC4WSiC+kDRdw+hVUWzMGQfAgMJ63ZuGfpBknioSyVVejTjlO++dR
TbDhffcoW4CMcO5Dv9K9H5vp/UYldnm0429lQfcP8+jsC3iZEE3AgCes2zXTRwxiVj3R72uuZ3VD
4KAi0ciSBxGDBaUkqj14+xrQDpGLN7xxaxNEw2/zCugw3EiZ1Q06bpaiBRzXdJGrB/WGtFokpgkH
LySg2rsDDbegu218f5Fe8YLxyhwJvOx2qz2rwm2yHmWGfMWgYSNJHaWmN/+ZzDsLwPwBeUUrXhjf
5PhHu8jr3cZP2tlviyFdi1gWV3ueYqe1a20I6NEkqMxBIXhWwLdTd43nVejO2e8nsRWJ9i0hMul3
Y1kMAnFS8wubo8cv1GwWJi17dfstzXGIav101QARV9/8Ae/QCDd8gm5Mo2BuuSXvI/8w2iJRoti6
V3vX6g1mfOnHakKVsxBYCUDjUsh18YTMKqRKTT7IdeGRCvwFUT+WEmISxzzYP2bBZkm/zkQXTN3m
12LH8Txec9/KIR6tNuNwQfVdtCJuxvN4MSslsOXh8yCxwJvHlIKSDuSvstAi31U04MK2fy43BRyr
DkXq2caTOiSeSmktKtyuxrb4UN4+DLFHqOO1Q2dLPiQlMrATVQ4SgSQYnHTEC5djNlxxeuRgrdeK
2U7V7CidBme/NOPRhVwajWOTVT0+uu6DYt57mifS4SDIRD6RdFrOiqETYXQTPH7QiZlC88up2pg/
uP15Z5816cNg4B664ncXnqVYqZT0Z05IS2VwMRMD9XA41VFjuPTH1HlJZ5Wy8iKiqnZLqLt+G5YL
kZRfHuHyysmC5RVCWK6qA0fpyQMFLIpUjQy/jBzdHN9hIsOMRn98Q/xLh8KoBr/7LyAfcTzsAnp2
aZiv6sODkle8FWPt1z6w0Fx5INoFG+JCIF97lQXN322Gx7Ig2BYDg/bXHpxwo6Hr+vuCNspJ5pQz
0G2GXmkjCk1dvltk5isnl/8EyMZeIoHaSiKubR028MXC0/BQ4l72gh/P+r8XC6tDGWaNzheymjzL
ZtkTc3iAE7uyY296jYmOAkm9mmnOLfS+n5sHw/9sryeAIO8Zmz9MZ8ktcJfTd8s5FEbc0m4DfoNM
/VQp7sFKCk9bRECzpKmxl8xH6HTXr6a1QOa1QsySm2n72dvC0zTfogOSBlpAh2ji8aUYYWZhNOIK
++9nU4/W6fE0c8kah2EMx/9nQguG38WMBZnW12G9KqJSHmU8ak/pY8IO+lvbSW+Tw06RVnMbmTVm
0RZCvi7qr5smertNMQ1gpVWgaA8pJazUsqDMNM6n9SIzEPkOEVH9boXhwnG5BkHSegjEBb+6qtU5
cHQDftTkdB0YmduyuqxQ00HZAGMwsciLKJYwXnuNLwalcgu+hKky0kiVed3aDEZmP1p2iywkUASv
IGN0U39oEKeSB4/ckFdZBQdUVbh7q+ojBzfHRNstqdIXFhU3dk5wI1nqIeApeGprCu440ddloNTe
gYZLPu/6KbbnS8F4e8wcGerKTphaW+c7AauCZJAIXD0NlVFqUzJcDM1APHnG1kwasKRppT326uSm
DWNtdP1PneJKK8hVE4dh/cisYeEJ/B8SfYNiOGUYxm72mxtFC14QsbFuiCc2e/Lf+EhtrHK0uDKb
Q+TqEY4ftRRRz3XsyTznIN/E9Pv3ftk/CsM5VMugFU2YnsQUO60FUWyl0fOKfwxs3FMZUdGgE+Cj
fMFgbqOhwiB2pEdjdaH2bBza4InuzwAMt62YoMxTVCaqey2KXDfvW26dYZ1z9baEDLA8GH+lRSQR
7eWyX8j2Zp97uDRKPDMntjW1RTGBJu76842l/7FNpsIjEXC1zLgC0zsLdepLeGhn0dK7vvTvh6k/
tUUr9E085xe8QwbEUs2uUFgxaajMAtkz2cWikn6ALR+TFFrZgftfVQDOVfTcuG/aUZimImYVoJS3
2qbAE5fHWlotv4UDCLn9OjBa8HC3mVE8G1IsXbk//oT8MW/HaFCTG/C6IGA9f92+z/mp79kQWBPW
Ker645FTAtyA8AZBbpuHrBUYRSs8DujTQxSV61dkEYKZDjGMxu79JYoOmvSOvxMZcGdopUMgWN3X
Z2mp9g/gYWxp6QTgwSXHWDsPrg3NbZJz3oz0BS4o6jWuzNXznEE6eD3N+Umv3fAxnMI3RlYgOgsw
y3Bvn+7Km0NCN2ipAbwmQycc/L0MhsEEmu7j9DsX2DC7E2zMazLw62uMOn0PkzGEiQings3nhsSX
v7r+UORkAI0b+q8111CLMDuW8nmRpupHadkLBLF/B3Hy4HsUhg+aaAm1B4vEx+1tGvfAmMJJ7tU/
+bl+IFr1kxQSrvyd0eji77ra3B+N6LY2krwnD9zqLmOqem0mvR/kfyLMhX6KbGdiqsp7Ojjv1VHh
u37fyTNcp4rXqgq9WZbNSpiU6bM5M8yEmiUebkh6o3s4/SHpKL0aET5HhaOhsNNM7Z5BkvS0WoE2
pkaI1GR4fU2TIXxNBJRPC4vPWsbXiMwHoaz70u7hhT4WC7Wmd4BoKYsxUMhMpx0u9xxJ62nmUvD4
qk33JF4RMA+DkJbPePgUCP9p4qTnVqJczhxXx/0mWgpZ0F7XY9QlnAIYzqKnnpPu3Y8rJxRPeeVy
a8Bg+6CU+Zpj6LUKGYluyHzCRxIq/Yk2Jv94mCrq6JuNlUUTOgJ+i71xGJ3pPHbjUwwHryPywpgO
/MTIiR0ieqCQDbznep/ip4ikNmt1kXeID3bTcIgazs668hPNk/sOHAkns5WyKD6ywZSiGE1Tm2Vi
Cxx3QkXupqqqs4mvUEJWPi2Z/Rbq6voX3+ZQ4QcYIOiNoD+FgyuPRUDpUovma7R9wsZFyhyc/1Is
j9O75W8aL41jNVnwCNyCSlZC4RMp1m/ZjBbdMIJ3MegmfPM/lNmTtFUMU8X1vhZWFZjYzXP+BVYb
5jCCMbh1qbBJcJV+/XHClDhHhkwij7IyNyaalkroL4c/MeiCNnmWIg7NxY2Jt8b+yunCKYHiS8VU
ydyb+Z9ViySqcM9ivZLUGs8b/TULVdlPv3E26OKSoZIIzqNhsG1BTjuj1eaGvGwre6pBLFv1i0NH
gwsW/V/Z8FidOkBjL6VilYvWKD32yQ3nx29OM1Mv9VCGRSKwqiem40cv7SEgMZ6hYcGeBis3F2nk
n+N6QOOKUVyNJb66QR5Z49SO5FkbQu3EFyanKcW1kKAlPw+R0ZKTtBXH73cWmpadUtrjGatS3RRb
WSVoh/RyXo4K6kgeFRHvpJDLJYGoVf7sGO6hB3n+0Xe8xkG8I+widPSdUFySr/Q6xPphqJoK82Ql
05Na1oEQSUHh9idwYt/GEzEfzS6A0dJyIPkqqqdAowy2Rbeoer8khaLw9UlF4vr0cVb5Uc4+hHpT
wX+r7UOaFNGQeNhkDoP9z4ltZiiUC/MUJFgJk/65k6K8hKY74vyPHMd66/Y5wwM0wMEbUFFoKaCZ
PnMQf8wo32rVJPNXdB7vtwimHmTfkojPtB+fDoBWW+Sp9J+ry0h+4BABq6Ctr0gnXUBZx8biqu5+
e4Owyy0sLZnQKJXSsLqVePQ9p3XwQ1/4cRo+yhVqTeYbAqgX5nnhHCkm6WbW8KWyqLr/2tIUdXCJ
vO5n3bmr82qK0cpxfG4MPulhrq3eyFfUfUL6doQc0XRpe+CooiBtNcnSDN9fgUfHeNgFwx75Z600
/QI55L/PbZ3QfbYnngfcEUkzikeVjGBaYQ0qjhDz+TC173guFXlHuW7H352DyORFSKZtxgobot15
JF1AiwaeQTaAZ62jLXXa+cGOB08fYOb+EnFuI4uibaFJkEf2z6JY/xD3TZ/N+kNNSPGdBwfp9I1v
zB3fiLmgMs4E2lz3SovbZ14z2OoKlyyq+nhNk6rMy8/FWuO8iCj7wUDTNcskxP5BGSVA+yMPzgOV
f79hyo52hcrkZyq2rlHhI831USLODRfwg9Yo4JPu5I/6+T6gBhe1OQaDW5pcQEW7vI83iFwBXGaV
YPQA0Gkqez889UoXRp84uZ2mAsjW4x5H6wwxa1d07BFrwQNcdIBckdfx2cDtsGfm48wZ8ti50zpw
O6A6CiSb/ho62WyJVxbcO8DkUiSzJs0IIdE7IDns7A8nVSUg/5qHuxyviJrTYi4QbL6QF/538tLF
HcOogPbYPiMA95+Aczqu1o9ndTiXuNna/JesRm+pvATyMeVJFOVMbLBzGRpUWaSRNCqc7gW/tKRU
aRHqQw+2xPsIOD4N3gII4mkgZ+mPFgrkj3LUd3GV5Q9z881YP42BaKn4bj7pLjzFwCAdeTeSeaTO
E6ghWaBT64wfuOQCX3utaJrqhb55BooPru/jFwHzF2CHT1XFRBz8aEwBBps2mH4FUjrmzzUvViE6
VYJ2p4t0wrRE/CqgY8+H2Mmsqy0ata1RhV+7rUBciTVpdZt2XgLDfPpGc3uHn3lbZnfhs/OF3WBs
wwVd2EBSF65xJDBtYPWgVcQnVFx6NpaUqEYjt9YTMzSJlVpFTrMn6Bjz7wGsNDrpOyA1bjTvdvIj
UoAw4kHvTraN9b5cfbOjOsbnmcdxi4zgjr6t0MygkXAU/VHk72PMaf1cK9jUgKUTD1IgbfHt8FXd
lI6GsHUDgQhA+aXrLwCIEmyK6U7LwysAed8CdKfJei91i+AfBqJIIcanW6DBVKGWZBCd/mdVQHfD
yNtS4S3dobSi1Zn7pVyM9r2SXLTQ7hiDkArsug9tryuEOQ6zZIO2R/fT0/ci+nrFZstNYVZA6q16
OMhiXVULVZilWIEa0V4CnsV2AtsPypblN2TClAhKNZnVW88PjqowGUWUL2y3mo63ctCXaFltNXOe
xJo19lTDATaTUYB1t11WLfRsWHAOxfinWb0TPCacb+6qjDjpfb2Cd1mvua9aMpOg+ncnwY2ce3UK
UeAR0zhOoy330ip2RlIwecJ0Pxl0NZ0ywuzCx9YZ/EoqlOXAyD5RZ/vXxHRPKHKsRCmztw+Fvd2f
veZ6w74Owof81CcOt8NAu6j/qJDx4WXZDfYfqMJc8jfjH35ipHcWjyhbnxrQRrAPxeq4JdhDsnYL
uG9GEeiI11GY197JofdEMWH/NJ/G79AK5lfnOZ5TnoB0swe1noiUHogNhhRN4wSa6bm5XL/jS46q
9SDB0tZBSKfvmKvLDV6hNdokX4ovMRaI2FLN40vzkCBYWw8R2ti3qComsaZvi93KzrQOhas7ebYx
BvG1DLgE4PB0pcXSdV1Gnwa8OBwfVBsOnxE7wewCFrFWVkggMJO/gGQJeWEm6P/DutFgEdBd3s28
mVy0lO5OxPmYwjgHJQizmbq7Owe6g2ZLiiHoOdsvEY/Ln1DYlpI9sMmHx1buwfzOGG3lrMUvfce3
qA82JBwEl+TJOxssYfceSw2wyLlchErPFYGUCHSkdAnsI4VyAbXa6Q3rWS9idZPm6fvGp2XUeQnW
yIkBX3J2u6+GvzWaTQqutDN5VlgXutk6mCqRiJj62WW48kV893R7SVZSDng2a0gnuEmJ5cpa0rp8
YyIEM25yyIr3w7iCEX/+J9F8ImcFjclLmtw9U4hARcgFLxHgNT8FnPcpWtXfH0+vhovxpOD4q3s5
Aqp6SBcm9+pWwcCTg8Ik6bb0YUdw0AIqW4iCAMMhm+nt7SfceV44JW6SWt/5CLdvtcWFuEF8NznH
M/vYUW6Q1cZdYMgzIVUxviRza4KBdt2/ODXelVoZ6ZURhcFRp7U15e4UmwxysohUTdU8gR6ZZQsQ
cW9ASl8DC552DDB56osyvRoAU44W91dcHQ5NpYbiC8cjd8hatQjTLbmzbFcPeG19hrJMY7+tjndw
Eoav9SGSKhuAbkdf0fI0kDM2wLCuUOPFGeqUD+4Zh/zF5cfN+69RwccZYDgGx7NOe6d3zr+S/ysR
3GuA5tKFeYHtdnzGdMiIN5GEP4VPppF7hLcjnfZXg3xZi7AKFgrdz4MqwIoLpy8UtJji89lrDhaj
HmO9lXAYJqX5QhhaieDJlgdkKJ72v8LjXCz2IR8TuYCld4w0NIFmFeF8caV1TardWElACiJJ1cxC
cK217ZjSf1mN5PvmNz1gfC4FIsDTBrxfGKTjD4H9So/wSpAoMo/gBZgylyswZOo8r8+pondvVKZD
ORdJ2Cbu6aZ/1Wogiwca7C4/LxiBlThx95mUsOoezrRwH7VU7qAWPsv857/gbPz6FDoihM1Tza86
TToRJEj2dotlJ0E8Z6T+lBUd6Q0stOWLAqNeCczWad4YNKz/de8G5zrFQ1G9SJ612UeoWj91HLb8
fg5mB9NwbakpivcFcCB4M1xanR6oTKDyxQINAdAGHkY4RFqLKmQaveorTgbWCm5c5BMeTYjL19y4
wbZ/P0MTtJMryYF6upmH1TqJKOonkaU2dkSscb/GevOc/el0WpxZvjCxoOJ41n/s8woUgS+AL6FA
1l3eyO572CXVbGm51U96rsJDRYdqSl6Zee0kBRo0rp4SRauBQLYZqosvAhda7n6FT5+BLPsMXhNF
Wl79W3xieiIg0DPohxVtwuV6kenUfT/20yNDm2LsjMOuQdlRnN4PNJKFy2F535etDp1FtoKNe6we
iDy0z8G9Wx3qxIbhfzoHOjfeWfbSbKdaZPxRCw9Wl/EodHIBC7f1zYKQ5plzSKGDn0azmnesqdSV
KOguEJp5bz4BjQ8+zkxfEJW+b326I/wb1wMnf4HPYhV3+wk8j9wbIhEK9Jwp4pjIQG/bM1iuoaHM
d7KjlbppwTVe9986fNFsjWtbZT+jFn/7nc/k24bkasaJSoQxuK9tQc97cuztiiybv7jb4g1tPGpF
rYUKTsmznPj4QAMz6cGT5D8MvDCBmpyz9S0ZDdCgIBLtKULmY9ZNO9UufK4dp1rbYfAZsVtNnru7
4JEspw7HiqSNZMYW3iqah9wVQrrJa16fLL77G2skA215MH9icK8B6M1al19teZNLs3M1uCENaS4B
LlfABCsKwJwmPjJxQxgvOLAXSH+XbPGuByJqeoiCK2a0n6vQh4CXnbnpGNmxEgsG5E1x/oSp4Ggs
V46o7RyjvFDKhCafTcj4UTASKjdWJ2LvJdirZwat17K6sIp9/b+uAJFYh8V9cyy3yKY0Bh9QWl6m
H7qC7Kgu+qs2i8vj0cpFuc0fInJ0XRg392dMnrWPSG8aVEG4DJEtbw4etDZo4lTWKAV576AZ8Gv2
yyaGrYDOR8PT+KrJFdJwLex3Q+3lMkDCqfM61lIzNnV8QEMSyDvJWjK3S+2VS/wx5Bh7XdmEStMY
r62KcUyVZVFvvvit96dxfD17l/99XJ9KpNTg3BlwzHbqUOFxlcqQ5f84faiP/8GOZfS6Ty3Jkrpj
wGP8+XxA/RKJp9Binvu0Pj1GuCSpLVz+ScFsUnGs8b4DKwhBahFqpPEXui36itxILSaYllvvOQwc
Pc5ivoGsr/a4KmY8DTPkM3NtQs9ezbFFevw/92Hxm8w2xp51b8LNTw6S5p5uCzQ6h1DAc2fp7FRR
Sb0hDoYMGq6oQakQwKYLpdeFJmjCFMpkY5XAluhbx2baFNBoNaIuxt/hd6f8hn89yF3n6Jdb7JA8
cjTIB1VddjOKnW0LyzUqR1wQ5eJfhPoQzEUT94lLTcKXqwrFbmnTwhiIj0YR2HKBaqin6L6u+N9w
qvwQisx/ZdGWujbjXeAsm7xzuwfeCoOzeDz7HKa33snTaFmHidoRMCyYNsElN8josGjuS30qBt2p
yxsqZaJmwmeKqJRNyXNkcE4yWewqRm1tQ8pHuMnsOSd1zGlBjLszA6Hy6BFRb1b6NJz9/x0tOFl2
0ShnoElIz3FJ8Gn+JOlgQ9Ac47ghIxYq09f4PK+uHN1iHbg2lA0SlRZiDZYFKNj6DrtrdN8WZT4V
t+VXsNXAJsWnRlm/cwb+n0hwAg8CppXIUMM2ULYAkYWdqFzvJ5UFWMu0GynQlRWHOO2SaZcAHzfn
USghE1+c9bNVv62VjU7LM5cmQ8wC8DRt2edYUodpODBsyomK8i9bSVYJDqbCSCj6iU9AWTowDiv7
6aTalFey/Jms5NQOTjk1e97IpR1q4Jv5QzGdgDelFqEQZAYeExXn9XSLnFaRX/+t9f9hKFvFzWST
tb3MGtYVihCB8t3gkdvUIDVf58+HBicU3cfjhkalg++VTS+DSBpf/ficUdsWyUs+G3hbKrae8e1x
YLQtQcF9q5UCg+MhOpNBU5qLIQZoMps+jjvdBBIt+ktkWfbMLHdceMNG6PODWqF0xtStqZ64mYJ3
9Pc6hH2Uy0mpCf7RC7OXoDrX6o80MaKa3CTgxHrNgIVABDH5SlD0xzfwW7dx6RjED+r01NdYayUw
ugsJrfhblO6LpYsAH3l7eXwPY8ZdJ+pCIXj2GMqnpxdQ22UyPYwlO/ruXnuyHSNXqZeNwvr3rFNE
dWCDuKNvcPRl91GwVnHRjWloB+bYdAzBTy9tofhzrS8iVpbauSv+hb74bE6tbt4FgH3oLg3TBZDL
Fm0J9s2hFoJmlINUh6Rczv0stNSg0Jype3eCg7PIJ2d9v6l42X5UMyE6KycRd6KhgMgZH9PS6OtV
Tz4rVAuOM2/FBh0ARyWevm0JrYWpdlOZoHBLY77WvWPUpnYdvmBmSxHCQ+oDTgQCwBe6q4iBV0Ib
CTOStAE8GNWDOD57IL0p9us3b0rOBwZ08cRdBjRaSDeuBgP3FoytpCPeZkCQx43T+YqdCIrouoP9
uL6BnIbN8uNYxpFXPVhkFO6JfH3FfyF/jz792KcHPbShpJPlqEGzItrfNHz8lnXDU5RrMbrJzPgt
tgEN/Rva9nrAq229N3j+G3G4Gu5mZu2FgFxcN5+j6zE8mezC/ixwuqlaPgH089FmeMx9EwmGE+Xj
DdZLOvUwqC1Vt5AK1fAbujLKB72kXljp5qK8yAxwWlex8PTqRRfhlXGkOVJvfLXXgClaVrZyWvOW
GxOItgQebDquSdoOPgQ0k7qne7dEP38qM65fRhCNbV0C1GtYazT8yRiFyjmmFtRV3NAVzYkoyTCI
NLtWUDvqp2dbxkFK3grXCveGjs/VmMYuq0Skj8bKMKOrut+i9/kD9bWbS/mjxyeIXMNYKD8aoRqZ
ueou5tWeCfv8eVWhYozCXuGtwct3HuExx4kZClDMkXifaiT/D8GbUBFxuGQU8p310FBWU/BASX8N
xEB8FoCGINNl0/c2xIHhAZofrvYycmWFXaL4xjsLVNXsv+6kiLO+cxM/8841caQZrB28eK5iLcuV
B1jkarjbTDT0fzj5IF1lT4WC6Xy3V19CcnUYgk092mIBENxU8tHZ7YcrbbatYt8ul9HtSgGzpuS7
toUttLbH81dRQaJCNyow8Jk80HOBHkGVSEYMV7MeL/ETrf0kPTfctrOmCTEiTPDQ1wudOagiMNNw
LoutbM1qD1B/sGlhMBRpEydd7hsP353dauBWb+BEUvShRvpkpG6z0Or+7PNe9OGhPEt8IDyAuz6m
i9vOxmn3njbdbMg63KiDNWLU8PbMN4tfRHzKXMmJaXh0s6BrvQOYzGDTgr4F8Aq4/WT8pB+qHJyS
tKKXbOJw9jDvgh5WgnpltXj1r+s0/d0ChyM3SEkx73IJQziAtpCVh4HQomJ+kQdxzHD8DLyhiiGx
IvKTqdgGaaUu4dl2xDe93fi/pXbIazFNdHLvYaWMMRFWFqDyasoxEGnDldPJTVi0TnmiAf80dN4l
ajyNc7WE3QxzI22dtuXZah/2xNYzQ+CXEAJWiltkHv7xjg5lSCPBjX+SLcafoFGeSy7I/mbwsABq
ptuk2YC/qui8dwXrJFGINuQnLonf7gKjzyHOniRZgv9PDDS+m0LaSDE+jyySrmODOjhRKd8+htVI
ZaqbxN5xh0EJvDjvQeN4ILEnv6X7zs/kz9sPEu2UiscsZwznRWNpUaoLNO1aIWAGw+9iua59Jdnu
8C7KCrxsRDz8kFXSLXJ0z++kMfuhG4fzIKV6+YMT2rM2sumWZamNFtcQkRGjMp9nWGs4UUQ2NVL6
imn9rXLy5B4/bw85jk2io8WRXZeeeUasTPqwR1zwCgCu/IWUN66pvlLEDewE5LIT5vBK4D4NzLgF
+cc8claEAWFrh6tRFJ469cTEdlUAscbEhxP8j/PsdXz6OoeneK1QA8jJAJRRUJqYjW9+HEZpWm+c
7Vf3Ln/UMbqkxg7Gcsp2SSa4Exs97cPV1eCnAFQCO1QrxCDMZVQKQYEz6wVd26HQWEZJjgYF2wHX
scJS6HMP6wp1Elm8OMWai/ZkVbvKBlVQOlA3+mGM9DplswOnZJUAb3aC7guteZmYne585KlQ4jzv
X+Uma1qaeWx51ypwQTG+mXEeiYQ+Da2BDCaI04aGG83FdE7uwaudbRPdq7F8RM4Etx+jrnukPgXg
G2zEYnWpPdkap3tZ4nszRscmBx6hTWlhYBOzUFH9C6gI48C2CVV0YXOotw9CAbrtPQEyzlD97wZs
D7uOhALmfqPUIp6Vu1CWV2qhgxzz8mAzKw8OTNNfnmhMydmnQvAIrZKSqndLAPnx7P1d1j6sdjiY
38Jmre1vclR7B2ZmPmwVQNTxPVwJYEJ/cOM/7ePRotffrmXDNp0fZHSsrHxGQFP46FB4HzNDWA9N
ACjYlWHiWIlsiBWAWG3X254FoEbeIQcYSzNJ9rKpFkpGU1uVOLVTjDEPzupn++MBi4dowKTQ8l3a
3mCnZ0/MwnhlKGvS9DuCxfRMzHkuZ4ANKn/iLNkVvmagLUEcFioW8stZeYq2/ELA1+2F4fYKTKoq
QAWxpyT+ngPDoNxKBSKka0IUrYsp2xpTvlUUcgFx1QuesJGHKmoc02DPDSlG1LMIw0wg1Rg10rkX
Nui/PpcKyFiB3rDDjhTlkHHchDuTKyaAYXjo4H8blgNF2mv12nSw2WdLcnREONPxE0QfAd4U9bZi
3g2lEL6uZ4o83Zpo43265NIvj9DkuSnweOyaDd7XJrBc9CGKurwI/9ZpEdpA8/S5J0/KkNLHG6o5
1NurKrIo3z6JStNo5sPpPug4fTRkrLLvYECGZHzAeib0HrGOQzw0FWaAeUlEjF1pw4HQvFh8D2/I
TpTCYAfDSbho/mJHLbVCMQQyTIzoM6ShfjFq2niX2e5wFA9sM3lyuk6TrVIN+lDum8GbZBOKadkD
qYyh3Dm8VuC0QY8Uq+zN4z9bqjFu39I6oneBIswJuTIPH9/Bb+2trRYUnjUHx62DgO+dqTmBo2dZ
dEUZl910pX+dUcDmpuN3jOIzoc4LKPLP/bjv/Mn+zPWSlDlGnloNCccZod8tErV57DC4qEtpsb/Y
nw+9i++VpEUnlnHwmFJSZeMuts7LkxXrmNuIAp6bj2WSR/XqcH9cRE3lGU6ZYjSrdIYaEITd7/do
bWg+TI284wncciwjFNlEbpLzgdKXYG94KkFgGCQ/K3vUF9kxlhg3KIRoTB85rnkJxXSUU/RHgmKA
LF5ewHgPb4pe6SUuSkdQckLMqgD8Pd+RGApOJi6geHX7BUmFT1nN1CIPdkgj1tD56mXi9QcgZzMy
LKBXeYch+jM2gDHmW8gVP7nL3F0+Qyfk22goCuPRDDrYKg+Bfkn8vvHejgu4/vqQGhmpjW3TVpEC
tCBU7l3uLYVWDcbTyaC+wQX6S9iITQWfhoi6Nu69jO1QBQh4sO9+h0XBPtc0Yn2ENS6dXGjRy0yd
cWk8dT5PZvuiiVyYaOGlf8pJFWWg2iDljJgfj66kflJf15ZAe1vTkipXEop7HD6Szt7razcX3EHK
uOLbYJaRytDSRisXKsdeuJpjMPsROYz+E0NA5EAemkfeRv36l0CvdSupBdywrASIDn21UvzR8m0I
jxUNyUpFo62asf6Z/+pptw5JfogbjJnITd1aZI+J8/NqnyyLQUuDG21jQnCPfAeqftIDN52YDvi4
LjZDEDsExD7xHG2tVKmwZofHzxp++cPS5Y4hS+TW94DsRFnBoZkTbXCwfm4f4Nv2BkrsTpZx5fUp
kU+l2cul3uVlZky7/g4e3L7SnjN3tZuhRbdkc/uMkjZZYoSV1fDslDum7CAabxpTB5sMDXNFN8Yg
ISQx/kLfEZOhbS8eLONPb48NO0nx8i79/e9W3W/Z69S2ThfUparNNfD7p/IzVkFrplz5KK+/E6oi
jq293euuVX6mSoWNI4pyWKzuAHm1Oi9t8ooKviGFY5VL13/KE5z8lw6c/VkpMUAhokwz/WLmc/BZ
hKk6te5qAeOeQq7WnLh8T2FtDsVjpjvfDtLUR0apRzHHHF/3y0L4ttGtjp22dnN45FRyHVKCJ+Vn
Zo4hCrptcJ4eoAyGymAF7pKUFvHXyR+Imql/RDuJ9m4msBO15+TNkTHLjXC58+Yu1jOOuOFG96HR
ngKdrPoOMk0tkpZBy+0VrH4b1LyUpybP0MgBrRFeJOzaIA1RiEsr1tx50kanBfiBnMiByx31Ttek
FpYmWjcCib5okecbFVOc94E1EOpvJFe5AmypAX6hoUUUVyStZbdcPH2h4uhuN2Xi1VYnpYUoS+m4
IQzpP+bPwA2MIvjFXkeOQlBNIrMXd34ouGtouz99Wx6tmlJ6bzpiZScP/44Ni+skKP5XsTOcY7qI
kuEqbmmAxAA/sQBaCPTAYJWSZyAsT0jVUIou9coV9yXduXrecKY7nvCWSmdYtvys4fPjRlM4TQIH
z9IbuzYFu/W5oEbev/Mja4fchj4/AmqoD0dgef42o7y8fAD5v3PafFO/k6BhXBn65iudqPlzIJFM
Y+7K4zUm7bNdett7LmqjP/JMCNx7WUu372FVg9Fas/ePgz0HueovMMSulmRRIWT6thfZkwmIidgT
yrrmoFcJedgDB4V1rCDRkHe4lCzCTjOGdYM/tFZOw0naBoxL+y7kXWibClIdyEmOE+gBQJd+hC+Y
ni71kO99AaE9qrPXxtdU1SDmeHZU+qM9y1rrD5zwaV3mau29t4ASNFdkl3xG4YL/aLGXS+W2wlmS
cUlqAA+BG51Vq1HWmyeZkLpO1UwGsY3K0HL7y4fKuLcykD6JYcjSQpWxtra1WdVEWlj0XszNaxvm
l1+kGT0SaShtEgwPrOis1503N6t8Ngp8Z+vszhj7bVgc0fw9ow54OY2hngTLEhTy+eAx9VFsxtsJ
hXy3ouUQgwDGzyQOw4OiqFQ5cHFz0Fm4bcL7DtDTViXTXUalNzpvNjKGX+uyfTjqY+wtVM4zP00l
j8TGHHfIsg8vpbgypXFhREAsqYyvUT3BZ4u1gKoyJBJu7z1EM2K6n2hPmREplo9KSMA4g6YtUCkP
UGonT51npHD7MwMu4hd1IEVOmKwKvtmxFz3nZEKgITJ886xVJtuNjOdXzGHSGhbUPxiK82YswrWm
lMXGKLgCcmBufnLNHGhB1oBz3bunOhuaMGe5oB6Gd7zMjEknpbTBEpaDAR3fHBT7mSsCv2+dmWhY
x6kRc3wMPC8efWijG5IhE1nCiWI1yAZMdWK8t1dBhmNxfozMTD9+fB2/xcRzA3BDFnLd0v9EgpD2
xAbAcijJllsJHWUzSsjlrLogkgD98wMUfN0OXMY40xZkYJHCDgKtBW1/8CQRQ1N6Ns7qKZ5aUXN7
x/+yAtCjdi9DGRPftB1EqRdwbtgEdLbdASqy6ANu80q8V9U7k3G68VbXg8aCWGD1H1kIMwYOTxiS
Bx5U+dv9b7E+NNuSbKoCBANy89d8XrUFLBh0+IikKQFmTG/xcJTOmF33laYXpRXwBAX1AYl+zpD8
VcIKwhpTzO6+PkfGkuKimk4XldG10g8niOux/fkv2a4K78P9UYjsu7zUWxB+vOKe/XqfIqIcwd64
weQK6la0cLpIsjvhXuVYmKOX7OKBVk/XM3YhezYcZJweMBJti3E06CnsCtPkqIJOGdY77v51oUaN
Oryspnkdasbi6LlzsARYfcGTPRz/fb8kagYY43vmhgj+Pw3521mmh8ZCru1k31YEH6UfTa68m8ED
qqLCzEQ8jOpBV++aA40VPMlvJKxeeDs6qJTTMbnQEsOO14nzzV7CRGzEeXfZ0QXnyKd1z/9giLFI
/OtB4EN9//HXL9tabCQtf1H2PEQF4OJiEYk6XJLFsZ9JsEAIfK7vx7DmI8ZxNIpYOYguibWAWQ7K
wN2dhqHgxQDo4jzD0YsbjszY3ZnKPZSk2JWZKwPGkJNVg4W5cSSQvbAM4NFrZLw/MYSf1IILVzmV
rRiY1pvUOlDxfFzgd08u0oQAnvU12ZlHx7lhdDXHdpmtMqM4ZGya3PGtmXL+9rtRL7I83ZvtsR7i
/LWQbLsH2MWAZefLLqakCVuCsBVGylNT546roQGUP/ABW8wunm5tRr40KAPGti+H0mx0ThxdWcK0
c1VD3YHva9mTkSycFBWKaXlfulyHFCOhl+2su9DrmyKqyCFkfQ8OvqPd+g52RtdEDkxFw0HB3pzu
qc+pVxhSwnD29iM+A3IZca0SIsMVQkDcXWEY87DVBpI6ekhzuWiSynL/cw2Jx1GbA7raedlaLdGT
DF9yAAqxlrXwiP3sOXbcz8WBd/bccT8xqrcz+Si7gHHU/SdGJHWMt9kRjTReI1OufyrTgPy0Vxnh
WuQWBETcw5atFfMT2Qr7pJcgXHRQAIxfn63dqWNmZPNDMt476n3VI+jVse3sJEK/NuZ1LW/IiaXy
VdfmpS1Atbw5fjn8OQs0pEqkbu1fDNcXjpoe8eI6HKHOTxT1RGoomjtVPhm0q3gXu6R5k4tJHAa6
+ubw3qzY8hM22JUGbhVkQ/2Ox9wa4bJrdqcmbcy0ohRYTXoaUjbsoJNbPj1IWKWCjp5Ddq9/Kehn
8t3aB1/R3xoHSLi9Izn6CR1jD7jdxdW5EvHxRHsU7q2JjfeG/4ffR2Yu1XvvoDL5ToAZd+OpLn+P
XeS20mp7wvDuHusq9+7C+ETa/v03tINnRLdK91ZzMIn0i+U6/vbRlTR0e9RSesoXrF9CX8339Ilt
QwuGsQVGH5Gd6vkzAyYkYtU/GF5AlnqRhKGAT2Np1yi8+pFD5R4URm/nXNTUEJBXtO9aWK4mpKbG
Zb55ayh+XtUNA6TURqZjNc0kbUZ/da50wcRscKlnoVQtyuqPCRInYDEsbn5sLT7kNIS1UWZT/HaW
odR8Lq4G6Shy44pAD3xog4O77L5gP5fJPd80ZfUIQcMNqb1XgXov8E7AQrjso5CPRRJhrjvMt/0j
c14IJS/4LWWmHC5Cgq/GtCX3aGjuIhAnPxAje2Lzt4CD+SJDjGCS6oQgbeMz5scdFiz8HLCXmEVi
aosKEncL9yBEHWiNMnSCn4s0sn3yPAPs/zCeylllt1qePhtsrBmfUOAz8Z5sDI96QJFqVyL+PRlk
fT56kuYdY7z7EUa9JXfpR5HVNSZ5bDEJ2d7GXIDJkHRftcNCtMLuGPx95TksU1qj/1p1/I0hS8vI
Ob/rUuEllQm2XSne8TffuUggEBdiB3DDDiqz+zOivnaq8zJi0DRvF9d3Aw5e0DtxhNxQu69Dcg/o
+A+FCtLv/aqvnlDKeZ53qNjuZWCulc+cXaDTSTO3/FI68FO4jM3Ewx2utpXoiDp9goyvhgFuIejV
CeGGn5bgiiqtjMWpnpoX49CAgSLKuzCi8XdNwbzd8Gi5pu5vIVUbQ7XQNmnu6qn84HLha3fLyRGx
sNHuhCFakXvgym3Y62PQ3OXO5KjCaiGwoQiETKM1UJPsWufaOSEkv3j8ExfBRR613ELx52GHvlN9
/dJsRpAY6hbpeoTM8JHpH5fYEhNT4tRbit2/VgpNreVb5EgqmUw/9k2Kqbw2NjElA6PgsI1eWSni
wfI+bV6gZKzxfgZluE0T6OUAOAHoPIV++cO2OB8AyN0KQCIQvWXGShRV2Ps+RON2+X3HMqN4y1di
kgjAFMpbpz5D/kgQnnmPCPsBH5z7taLOXIolUlfNGh97hFIqL2JUwTm8krxQWcWJdk4wiz6juOJQ
E/mPRZa0XKNj3M5HoCLCqrI7jKe+ZRGBpxuTzoc8Hx+MNIauMINEJ/YE7Lr4j3+i/S61yvhIuAwX
wz4uCzgVxIGWckl2yVbLBDlFiNdXyDM7agvJqJZ5tkeyPXk2xt4ODTrEk/q+TzB3v8VpBUVU0FJR
Eckp8h16YqlueSThDBCVWbnW6761KzyxflscWAZ+XMfDOrlQSaQzpsEG7Ln4cq8TfrBVxg3R9JWJ
MFc+WXeTUXTEFdhYEBrza6L2mbbn3iglFKwKM8at8ZOpNZoKYzs/81nS1e7LFMKmQcvZBw/gLODR
+Qm0OtS6AL1oaR9yrncPqym+X+S2Hpy2XxMvfx2IXPGP5+549KK2+ewe9c5L5RJXMQT+u0esuQPg
XuHqTextVZ+WIWjMd3X6n2JiycHIaTmaNmWxfs8D4CYoTvVr41VEW6kvy95pnelnna/NIZT0UnIM
j/jzGaViQmokK6OHq7khBN7vRXMwF4Al674vMSQfCSzvS78BihKOUP8Ps7S/AB1o1+yMdJXueR4h
Qad7h8pYPIxCGn0ww7PQ1pxDazHX919pjy2SWk3mriIvRIvtVBDGc9z+sIyn19QpAyW365JeDMLG
/fiUwxoJij71sx1oJO8jNlPzRXiKxz1fsBMMkBrTUhcxveJsnbGh7dCPPKHvWI8EoHalCrSad7B2
qP2crpI22+KEgjkSrEGDC+De5N9k8DmSexqBcPzvZglKWbHFkn24EqizMWpUisVnBPFYbuJqzVzS
uRNrWVK6spBdb9gT/2ICUAAxMXhk5UPr3PEEFLx+BUGrs/hbsu4n+EohVkquvIw4utVSsJYNg/nA
+KjoFdn5IU2uUbEupf3X6Eh/HpUIDR/JT4T+GNY+xYYtEoXx7o5e5J/12WQTuPg+ACZDPhEEokBB
HZq1MX1re6EBrB6oI0RR3HmUp+K0mS5nZ49va/PlO/cSXBczEgBE0pqFcYsZVQHdFJ4FpLjbhNPK
msMR+1fMGTGhrSpaxyAt4Q18TfkWtv0AhrhZ7ruv28/CbyqTonl+kr6N60EL5EGtDEUde/WQCO8L
AHPd3EUjzXFPk4KcDx6gvQYjxXltglHCBuEly02Bsxk/BEMRQ+aP0unpDvLrsutf5++aPW8WGkOF
xlIN9HWJyJdJVo/BfME8QhrA0xppxfqlnxnLYgQQrKawTWCUVfbab08qI3dIQZoMDAyZbzE2BmAl
eMcdAjunW1uKfk9b2K3Wdj6ofBdcLhL8ckFtpYOVrqjDf9sGginnHclUrkPVY07r6UNs3PyuHt/Z
bT+/+ydf8npvV0SwhUsc5OZGKIJDlEcXiqrz63YjuTe600cMyhmeGtS8WntfyDWUOK4M7yh+bK+K
IcLP/gszsSodQCXLHCgayfdAAC+FEH67LkZaCzuFXZ6DAdgwgRaxdLL3Dup7dubInxv9D6OPGnnV
rMWFbzQWU7HlKWq54kj2TIh0ySIK1mwyuqt9+IZWUvGWrN0Fef9O8mLD3Z/wnLMcx1ZUkiLUf80B
qsM+KKzUKIY7fSnsMiS4l4NqFVcod3j/INUR4LOhpknw62BeeB9IuBqMwdOPUpTXRMfVR2/eBfYc
DFRCoACzlgV5fSr4+BzcaNOOkE+2R9t4To/gY+5W3Cc3K+LKQZ4FjIQLhd2RFhnk4PaAUO8/mKnT
AR8msKua+So5Vef+wv7oeHq4H/Apjy846BPIp5hu+7Ke93Zmq6TAAOkEUu3o69jWrm3Vja3ytjcW
vc9oLEIyjlkUVKh+bB1J/00Vug8SJthl54w92Y7uQkA+NAt24hqf/RJF0maZo8FIQFDPC/BuRs4V
UvnapYa0zd9QMUhGpqx6TlIX/IFkCsY1s3DonG6CQ/0AVvBv3IkDElvdimm9A4aZLneB+N4vtll6
lgcsanDTBsyua+6iMRJXvO7mnIpabkn35PzEyc/EtTsWPeKUf5XMoxGP2rvjN3ntF1Cs5UGwVvPA
Hpj6J97wZLmqTzV76njQST9+/3n3I1XL/CORSd5bEheg5c0ssN4bzIjb/7Ni5lrdV828vTsyBaU/
svDJfaw54r1F5ecsZDe2WgZe7oDpsPGhhmYwLoOuQI1j7yJ1yidw7Yq+G5S6ZhEVHK6nlwIxr1jD
RixOVO4zPciaP70138Pulv3t2HJftYnYocnprhYa87ysh4s1KbIEPhvOK0fXVer+VJaxNqkSQgkd
4Zh+Gsi6H4GlFMgCkBummxqWNP9KfSk37+lBPMysAqhJ4H4x4V+7U0rGpH/8PZSA0nsQUBHE883h
cqdWi6Snh78LHD4BJkQGMxgk0WYfCaYuTO+WeuNo1oTZbOh+7IgRNQpimHLzZqnqi2qvQCK4Qi7/
XCZ49Tf9oGlLTiEpOXHzv89yzze4bzL6+lEKPQrvyfSPsqVSdOQkN03m1+RN1uewl7Oyiqa8eTra
iu8SYkON/YLDtSiJXva1FAccaZelMMDUYCr02ug6vv/Yrbf1qDIuDolcOtxHp/9PJGJJqeB9dJhi
O3O5XLGRGK26QQdlSCAd4ILs2imCUIdEWJNHqp+miV5HXjyvHvHOC+XoKS2zJZQH03NQcGlzSzxm
/9NyWcNp6082ZWRMhPv1RlyUNf5Qzb8+b4H3OBLAuMl4v91u82ezJjzhDUKxf0w96aj+aM4Iad+N
dWsfer6ASP0mvNRmTMe9VUqNBrOqK948RDFabtIMvhUyABRVelHeiEQviA+bjNWjWhjUxmaWrxZn
NzoEXebZ8w2/+0qsMUzXNieIkbb8RovqyXudSjQpcPVFIMf2buM5M+imx8qArMgHQapSzEo8jWPM
76AICNjZM1pGA2Cm8JO5CCOkKUCDdRUFrcvs+hemuAPwNENIb3C422SHTcLYlFlOnT7wSf+GjTvD
wyL3MKL3AxXp87VDOdiWFTQZfkeR+yA6SJsQniI8Nq6FiVGVyAqo4JPzZGO/ZaPNTZwiJJASJPos
YShc0ahZXg4IiEX0sTe1OdQoS0KqogJL8EVjJSuhBIkzG+b27+mVEBC9dREi8Dx31rLlT42/6kSI
3U/3aN/tSqGv/Fcp3lDbLgSj/ETXXBbJnAGjSLZA8PDZRpQCTjFkv5MgaqisZyZwWPK5RqomrHYY
oZMvA8D9p/a2mKL6pBaY+hVdzu49uS91fr02YTJ9ucB0GWBq9TWzdafsjjrQG8kLGpuvGPdAFbiG
yfDL8g0ZI4BTNtFHEh771dYkmMI4qLRBCyINux/ms77KJDOTxqKe4XOOwml/BPQu7PtMXOsHMjem
d6JYMzml1IfXZRVrqSHJ8ZIC3lspStfeuBfpmvYt9W36gSfWTH+gP2fB3L1wL22jx2r4F5QLKHbo
48U5T6cg3jxWkxy8MNTijhJSCfGiPY4QsUAiU7nJYp1FMALOY42an7wczFKUyFB2JhxJHPayTM2Q
OjgT+4P9fFXTq84CTaCHz3fblM5t3uJOhBSNrubm6p/m+ItkOY2yf1yOUO+uRbkU9+hTa2TF+XUZ
rxoaKZDfIUhVA0xbas0znWTpJNkPE2ac6FzfQhMbZ6hR6jlolOMw//jW51XP0pTgNzSR/d26OFUC
qFNhq3oPM/OSksMfYApEfez21Ox07KN1cJs1P7o8UDbNge8UVMTmzTqNKbMQAIHnsJVrgXumOVGQ
M70aYBxPvIlm/L5JkXRaF8YoIMiCGAxEZVBnJxPz/3F7cZAxNS/3FQhHcSnR24nF8NBHgrIG2xzX
1uASaFppBUPIRN3zd0VlafO7dRcjJ+pQ3TWlVywz/tHljQrrt1yun25W82aTzsBUTuaQXR+/ckpn
4d6eQlFQlDwfPxkxEMmhvlOceZUROyLFs9MoAdkeIUfZ36lDG2HAN4AesciUB+z9GcSMNr333wRX
ZfsgmaULRD/ZWQ9iAMySY22ffml6b5x+IkM1SHGO75tv0GjzUSgeiLFUGdvblEK1m4kOqKosHquD
9oxxVi2Pm3Pa+CwW6NZJEok4sk7JJnoaj37dfAmex/6+bYOhXAOVn9SmqaOONpdwDcV1AuVsHm/u
mJf/k47RhdNHrs5vz7ea5fzcLjGi5EQWm7hjRZ6fgzUfSCDJAhDuRPHcXMbk8TeuiZO7U64JJdJQ
QlgrsC7kMcZ8Q34FXLucZoEX9CZJk4z+52qR29zk/GUBPGwhVU/+2jdf67iJngwZCpI5OUVAHjSC
8rLJvQFt5rH0joGrFn1KKoBq/4WwlK8XkFJ9staBD6YUXktypKq+x0lMBQN8bEc+LpV2YYx1S4nb
YzRJ5YPjHXUPCmoNgoi+szLpFZbJpeucoKvhAbQijvdvG6cNnrvorL2mTeDYfl8WN/OlR7mycU1F
eH9rOo/rlPtlz4mON2LEfjNOn5/bRcThxbeZlutftjZSKa1JqYFQe3x8Ee2LQFs7ywg1U7PB0KEq
Tok3TtMtMyNfacabNWjWrECrCOgfWUzsdvzWtpHtQJ2KhnhKHDhC6xOhaaZQErwgV/arCr2oG4jn
vCLJZAXZ3llshTteI9t9VOlsEIS8easeDdmxmwRXM5m4fEcPHa0EmwnayvT6fTi4aJ/eeTKdKYbB
QXJGOkr5pvLd74FhR8ubw0QUwlHI3jrGDvofEEH7TJ/vNZuG1RfbhhKN5G/Lhrrb1Bjd0dVVGSXv
FpMx4taATA19j1vEKd8ZkyHuJAzrR7Rky4mZUvDbGievvPWwHv+w02Z/cmXcMytjpc2nTT9p4PJL
Sejgo/n6Q8l7cOHsrIVnoPxAl94gqLfp/IAG2dNWidbsCmJsWPgdHDvGnZcx0U10TYcFTBWcs+JS
wTq8PN4MWKO7brX+w8oQk5WyewN7DeI4ZrFxW2fjtsnXi+Uwjr3Xl/7Q5unmtg9efUw7jmZpDE4C
SsEsk9s3MPY4xcl7OAZXYp/gdSG8jYUIHFDD7wHQcyDOtPiEl8GU3yp1sULBJ8wRY95leMnbTvlK
OvEiZ80goEt+TCC2BI2mdxPzIRC817BAytzYbbKVSJzvqPcJvLR0L/H/4ibRjMLjtvKprkFnTqmW
OvbzLZOfJCSJYbaWDWhzey9KeUPwZ+9I2D0dtrCZgjizP5YN6uiwdiIWpcPbW0fnUx3ILP5l7OZv
x+N1U7vXuITO+24Qe/+h25AA9WHGwDOqATChAhB4+mJaWC2h7aDHmviE0vj2G3IkVVAzigRxD+LT
uChSoxlzKn2juU3Q0ACUiWS+Em/p5lO/P26a/x8eCDp19EUpxyGtXvAH6EYyTa58W0AbPtYPyR3V
XZDMO+xUQnnF1+1ubA2V1hCYeatj6ATXe8pI3kEJJq/eRGRsiDhjPzEZVyNxujoGuiBxmnYmg0xm
Ll3LTD1j5/FcdG8vqxT4VDzWSmguLS1OG0uKcW6S7Qhj6VctaXZ2z8IAnFVVkufV0E5TIP9gTG+s
pJUe/Dei/K/qx2RSoMlIphjaM4bLNx7fGI54JJpkHrmzoh6Q7PRMwKmnDxgqywf9NhvswWgvtgXG
2EuwNANqaVaIEd9kRl919G4xT16xdLsFl5R5gk611fY7lMwAGzTNyBmzTUyQpRR6+0sJJxrqOYjM
F5INeulZIm9gx6405HW1VC4Oe809nmFKGK1nSVy1GsXOXQW4H9/3YuBPXX9K8a7Ab473Ocr4Q3yo
UQUSXgbG9+vpQgEBs7GdF7AA1+k0to2HfGSvwMBMgwjBTzeUcLH2xVeUy9Iq4gsn5ZRKYYF/X6a+
9YqWbwdj4Ks1b1vBTiffcxGY396oQ4uxPNNYxby6/za5GGl8nfHn4s/IL1wm4r3nNUMrSFIRr604
F+HbxeHM6tLPpRxkbzrDgUK54KdHkUZOFjBr6v4DNtmndKgrmCwSCmE3MClywwuj30XmV/TgTyO4
YsoToRgzmiQxs2w/F5STxndncET5qoFkYGBzh54HfN38cy7BnAIlkL5ouOpjp4MyH9qsf2MDso1j
d6ZRmIPru0q4VG0LgSp24Ftmp0ANKwPDUXYZQYYbQYmLzSvs5hbHz0EMQRy86n8Ty4xl9liKWTu6
RC5/HtPAUMhBDmz2HCKoB2rIXabiSXuy6E/rZvQQuxwEcKZb/FmugiREx9KdCK9Wm1Qy+5eCzZ5j
Hmji/LiKwOvtriYd5F+TOU/iblC8EgXpyivyAi6pIh9Z5TnwnnXwi7MBtq0Zedz8HUOChUgI7Jvj
85HCiRtjXi8hPYfuCB+G/6E40M56kGpuBAzyt/p49uHuRy48gjiqSBVWh/OyyYTLBZ6m6sgZwaep
xMh9T9impaJGraPNeO9SIh7OxgfKeMGobcAWdhs0sBlNd41bfok72Gndaj479H8d0+VvjJjQuEaa
obnfETZvu7GEp1O35AxP+Cs5xrhDXPWlDcO4cmFv4zdr2kFyuovHW2CLKF6NtRafHBLtR8LTLX6D
pBMhH3jgrTYxuDnhrELZw3j5VADJ+VhRFXQyaA36hm5x6k3iMchib1x4JLtQZQZUoRVGxh8HQCYb
tDbOIctTP59gJUK6ZspSOghHjCq4TodeyTr7l8S6LHNFCuFzkCaGQnKi56B6jaQWNtw2LBuEbQd/
PLc0iv3lgXPvfca8HWkc4ufNOvs7cL55GNvOUd2XV3AN9O4UmOYQ3s3Xfm0Y7VU23AmOmgaD5XwJ
X4k2mMmYuEexsu6rK872T4Enjk1IpzLhEtCRlnk1IFbmfEWpSqbvNQwODM1ZTzCweIAJAgEv1xC1
5vNABjkBhM+S0oGU0dImHudX2qerWkSWhKxGpJ9bGgTCd3LQRF0abBds2IT22yP5zC7MGAHmY9Eo
5gfTmx/BXwHG9A/bMpP3YDfPAqfJov05xYtcvNbA40QChEjT0GlyPAtflBhI4MlMuorS5uNjRmQs
z1HQk6kwqTqMkAVH7BKS+qltIRAjuAreNnMfkjvMWNxPrZxWXTsr90OhKPVxZq8G6OKy0bhREjfS
H4eHN2Sx5ZB9w6ybj+9FBh7QBWOzx/158tQJd6LI16dmT8ujgMMfbEhNV6O+UuWMSLwD5JoLJ+Nw
FEYPobWSiQ3hGKxaqwoK9X9F9l8p5e2ZYfvXVavKa8Rxo9xuGsgo7HHWpvUI10pPezFeY94+Y5VS
yb4NomcTwEfLljWf4PrqNUzfQskNcfqHoCniaBoHA6jaKfYdoHVtdWZ8uDjLOjp2dLXJBQL20B7T
herDWA22m7JmbFXB/W35iOnscYq0CPMg1X5UGoMCHLql09cffR/QrpVx/36TpsRvqXdirSqSvdDU
pPOT3qcpk5HthnDiK28s9EqjNOQf4Eh5dvhGgHiJR7BMvMgQgFDN/EiAiLH4cquEiNPpqCCwU3y7
s5fGDi9cPOr0K6YpXIHrNhle4H2/5gPrLIyscCW12mQJ3miA9EkHcAQrxEPsOzEe2AvzmIE8wMpF
ZNOL6jJNVGOEwooz4iLwcclfJt1gG7CN0Av51BuVKGI0r+HdMq8LoAF/9PzOpN9s3hqjg+uDHOo7
gRhTvzqztu8C42sMUTiNm8HGydTVhKQT+46GuFdAZ3KYsttwdQgSq/epU7L54c0UGZ23ztT3dD9K
k7WrimCWwAx3tF2fkhuxFh/GwL2lZSDRkKbPnX+NqNvRD00uU+OGlaPdfDsNsNaf2BTWXRCuEmaA
CoREJx4sEC5nNhr2m6T5nSoYYbRepTwcaPhcjaDrk3hrBncEiAErHDROyqxuWtvIpi50TVFkHTnY
sQi2hN5JJU69uu4OZH3sl5pX9+0WoEv7wO5S7N+vjoHtyJvwYtztoqGPmWVKg/4W0KzDXHPaX4+8
SThBKMt7Av+/6QHs+0gFjqfovR1XqTtlvzufdFojmF779dKMPoFSQT3lLNLczc4hfIu2886/AlfT
bogfIe20IpaZVgeqBu/a/F96IHzyuTKhCtChksY4qpHimvkzgXsQVREj6gD8/ns1EKBI9KO+Mu3/
XFvEShLSTuu7oqT035YWvAAelpfZevDS+o5Sz3mX0XMXClRBn2VydKX3CFi8QOkUyVif/2qTo+uJ
2VAkS43KWym9r4GYCralU9RCygEOuwJ0OESlg9kssPFTQ79UimkZTUShUDOnpIeLrdsKF5by2a2k
qfQPAS1rjorCgyXpYnqFWMgfkzDolcHlRfRObGq6n/I0+4nOkuh/SDpa6w2C9kNGDbzbr+U6QZbH
631ELLDQb2lx23m+FfMHfGnuXiTJlQ9pbXAG1DGL1GaIn5QjMEsyyFzUemcl0nsP2430KdPZOGKr
hunkOryBNK4/dN39jFt+67jH3mijjKUy7VWAazLeYGtKNnjzAtpO+4F8sMUzfPMoq3oB73J04qF1
mYabJrx7L4K6TYnKs6g57WZ3/+CXWitMCXcyOC/NgHGheQI9LaiIpHDr0tB4AF7zhsf3iRUbHw8J
IQpzaRlMsG2b6U0UuHyhmCqFhnnB3S/DSf/gGaKU5JkoaQ2xXN5Y51sSg6yrXtfJHIZUXuQBotvd
2e0p/+n9P3Wvu0UhD1YQigT88Uu5YyRVSOSfof33bmTPjdHQ/JJk+9TNEhyXpzyTJ3KdyKYg16z/
7GxRPwoXMyHds3dE/1LH4byfaakoyDHSXdi50lw1onG8mVgFa1RsureDjpc1QssDxzOB53NQzoCJ
h0FFJHj+MpfxA2QqWd/0DMf4cNiHVirOgFZCRlQnsByA8aXYQygnolP/6j9+VHHBd8aYJ9unM60V
FyPjFQurasz2Fc1X2iSIQhALPDGIymUrCDUkGGDPO8Pf0rCk+VrNC3NRhq05SchUUaF/m+pLhDob
/lduATABAj6UvP8hU+1lya8jxfw/0YjJwkSzT+IvffJ5i6Qx7S9MrOP5iROkdHft/jFdmTbm8gye
rzFk+8CNPDqT0eTKz54zPr1YIJFUzDS8EBzp52H580iKD5OU6IbbQTKKx8IOmA4UIusxrnYnmHgA
6ZHMpEr7A7qN4z44DtpWuxH/cQPjDGjduOhLWBdH29e5lgDrEvgh10yjpjKcTobjfrZBGVRMe1IZ
JQXoQ1unxWUvbv2c3FD7iLB+zix3m9lbROpsM65ITU4ygGEtAHRGJygZZdab+8lkD4pTCkmE2v+c
c5E6VPnwHW5DqvnZb96E0g63EPqyeNmFJBFIyY9cZQcrjq4c4Bi8KggUzrVwjooql1pgJj7FUV2X
kTmi78mUNG9Q6p7KVe8azbCbCIIxcZMUWUURw/YG77K+NhmoSbbg1fVWbsWXbUufuLjAyumJHT3Y
doUC+8lZrfUYKiFaX/6vZkAvfVaX0Tf4Rsw6CANwSZHX6JgzcuklYwMtRlO78NF0vsQe8jNyXh+s
+22sulCfWqNzVnnIXX+aNLJDffMASB9NMaHyJ3RFnNGC1locwG4wWSOnTbyxXT5FjMjob9k3vX5P
xzTMwJ/j817ssdEJfjfidujRPoqT2VZIztRZLHKRYl8MfPBikXl7GPKhOkTVWpQbsWWmD/zg4rnC
j8GQX1NCeNfVwrg5rK6IyIb+lki3Tv0RVsHfZac1UUdHf5xs3NEb4tQ+GNPuoiK5YBMubKzrmDdy
9CFgRrM4pldhuRuv3E4G3lyje/HyNBaJqE2Pqv4hAdXQYDmbSRWyRUOIdhZiE6MSEbZYHMTi0A02
sONPF/TDGpbs4EFJivNpvTNYJdfLSUS2akF08kPh8KdYTj0CeJP7ph+HWHMbeYSkGY2nIK4O3zBQ
8M0y9LfuWEEZZq6SXv6370YKbjsq6Dg3NJCdtIkAcqIsJ3Xahss4LBYwL9Vvp5XCOpcKfCSP8hWr
lNFz4/8kSaH4rPwQymDp5yrmgXhMDARMHkf0PsRGYQmuaZb5uAO/Ubu3gJRCzuA3Cl5ZPjxG6nJW
ioC2duRnAoNsGkxy/Okutfkpz7QXU5XJ25IsxH6dY+LF9hCFEKggWYVYQVgb2XmQpF/qA2j+bLvZ
cq5sklSjWSiMSt9H3b1EQnyx3lkJFNpNzVT5FjZ69tlDep9Epu044ENuHjO0LQZFP/Uhl1lwEZGh
/q/QVe+bS4sUYxgc9YfALeDT0jP3HtQdrkALwXfYTUkOjJFmGHYOQrWJQriKtDVJLw4ZILM/3XfH
Q7XuOY0O9cM6HIEGt3R1l4MrqLeGln1YLwZwFH68fGZhNwIUA0n3jga/rNOwOdVjaniLPX9ld6CC
zrM9Y9PmxcpsIO9KWBhYhUtDik9ZH2Q0AmDY10WZVeMoMJs+Nhi0tz85bQ0P2s+3OSlZhDLUKOUZ
M8jx6wCXl7yJ4guDa5SiSnPUkqhwqR4N6vbToPYqv7PULKGBUvoJQY4/3DvzRDMK1Gx7wZcRXESi
1VSS6PguZrTNd8obfWONwHe3fyibSfOtIp1jCkQ6kSp0T9XBjm5FH2808hsNAXTfAhn7adL4Yh+w
DzbVDpQKZHeM0Oo433oIDJHM5mLcCWJ8NTUQHImJq1YmU6Iwr3XwI1HR8Die+9fSFwHr9moImMDs
DPOrmulX32b6MRJ9aMFJHqijrRnfSHgdvc6++95YpCqPqVM4b5x3wqvqHK6D7ABu+HBFXdQdRBSm
eB7+Fw9v+UXWNK54spxafItXfKD4R/Y7DvkGaMiNgPROJPTqMEo+CLrXXvQ/M3iwKFNOS+Tng7Jy
rJjNUrkkaoRg0AOVYxE8/uscd/S3L3ABfZCkU11lO9mPG3+DDQ13xTjLahesp7j8cUiAzpxAvxfC
ahJ6ACcc8V7MtORgPuo1HQ+YRSEcuw9+Kq1dwkLE3bqsBUXjvR04FfjZ54oqw8PDBOE6M47kYCLn
PjDo5EjXwRe8hqP+VUtxEGa+HP1+6QC8xzOom2u9p1ptXDRwd7g2mufg2eWkzJZxykm4aUByea3F
DoZx1FbVYItPLJgC74UhK1T7GDneUDkjP3eqJMGa5JtctcB1H89VBratunHtPb1be+mQQ3mxMV7Q
IoSFPXKdkhBCHxLvBJu9bwjgzZPf4Kq4ws23Ar+XMjYJv25sedmWn+SvePpuC/z8j9FaDmcOjlzs
6JfaxipYIqLGH7z39FvB5i/bIs+m0Ys/n2YbYpHbbzqY6R8kQR7RhEo26xUVwVcfoQbUD90xUtrR
sOzxsF8lHtYglTm0R7A9t427JDPC+VCj1mWcm1Suf6xnYhdEG0AK1m0dTOUzjFl81LG/olJC52z6
qYOvuDdfHlyCKLnIACG/RAl+o6kioh090JYM4kkMpEncyZ717DPg2Gt7bLwi9ynvMz9YgraZ/FlQ
GHQhopQQTp0/k33K0NM6N03wiQYn4fNcy11yXDvSfWFr95BnwRmitC0iUn0LHuaiGaxGIH7mV4Fd
YpbvvSV0uSfeWGVexsgdnQgKoPEqBqsBXO7QgC4tiSzRVXIjtR91SRyGqOel1VUOZccTnzNlXJt4
OyQUnTHOYJZhqCxyDdEkA/IM9ZIH6NqMbwu7WSJL3wSN7cs7Yg6GY720t+H3VcFDSYi/KNK6XARt
ernUZFHTFyfFJaT8BqC/FmP0NP+ZgpGGJJURh1DBgB8moWDZsPRbe/jpzuZc5ufmZxCH5rkEl40Y
fc8psKvDMMNxTPAZCos9q6m6AuqqsY/b7lEbaA0tNRwaFW1KqXp26zLeew2qdH9qJJSo7DNNSFvW
fGTMK27j28fUWo1vxZsSLBUefIBnKi7QbOXv4hWiauvzFNv6nM0xXaKFMD/tGGfsEgk8myX0K8i2
aSbvZLadtk0qcow/zNJLCqfUzbHWmRxShvJnJXMxBryWmQd1r+qzhENMlmzlLF9inRF2tMh6Ikja
lDXL3MLD3oGB9VY2NnOEXjaop284v+jRQBRaFmSYSqMXtqM7XGMFsQ2i+LI9YvHa2Ro547kqqoFC
3NDo7voBVLxrYUjKT+OMywf2FbkRy40fbQRHS50rAv2XdhCF+ogwLDIQrxs3n/n7F6N0yTFbzxn4
jaA30cFP/AVI+Aq8beslU2leSTL8S9uIEvd7bYhJZD6aXbyLnV/SnVvcQlrmXeNZ8ONBTwYG6VAg
uacyKslsXfU6WDAYMijCHnrpBRVCPuaxNvyrmH9fMeN3YjE1uOg/zxAsaKr2H+1tgWEGCJfxg97H
+kSQnLDFqHzkal1ZdbMJg/6EhGRWW5Te9VUJpWypZ2D5sm7Zlzgz6hurlJ1HRaBgI6TENOxwC8vf
8d3yGUHrOAckAtYK2OizAjgfIVHHOXVcm3dNEwCMNM0GmMZVRKX45jonSLxbdUtObpbNKPPNVnPQ
dTut7pA4LLapWd9Zb6lIVX5tdlTKDvg3oPVl6HQa+OFrzjVieW/7yX3nu1P1FWggueu+7knvvi1Y
bmGLFbBYr41WyUdnk/3zMiUl5m2lbYhLx9v5OUY9MfT2bJMdurv5hXJg8eJ74HkWIb+8tKHNrTlt
TJnhwUoLUtHX21nLzW+sLt07fR6nPvwymPuwdezxyfsKtNZH8kGNe25Qedhy2KPeKUWYwGSh2eDE
QsbaP+PNbJlBDh6/kkUG/gP9Bt6/POL/2eh1Tm9Te1tTXoo7Vpnk3YeyvrQxrX+9kPaNivbdbWCu
9tW/TO/ZXybbFp6cmz3nyHGw6p2DmSX0gui8B2x9hT+QA4UvAK+/4ivDL/kdBDmpRFYzHhQ1Ev8K
eSvFGBjdj4NoIKKkl7w6OyayZtO+WWD6tVaWyFvbMqbcARASCDyiJZwFJVvMnp1mEDd11/+4W6dP
MyLMaXy5+jaoeK4Wd+oi+CYoS31PmlYlLOiC63ZAwdH1Jh0QSaJ3XT1dfsUVCKrE48XML9z2Aywb
RLPS6flvnpTqdoMpuyU9bHJfU4DXsOJMxb0MmB1wjc1nqRNToFhR0wc9MyuS6eaEBM//HgjHVcDy
Lvbrgq7tMDNbB4plu138Ye8R/x4EbMpUhHP5ZusMNtUBidy0UHCpl14yqccUcb428//4ziogVeqv
DOLDcfMy5AF2+jXogHr8O5+vEn5k1fY07KVWuQ4bM+w7nTb4UXXiMWt3S3aX3COsZYtO3sTPxG7p
hBVU9UWg1RExkykcSNlZmURKzCM7A4mAvVywgsOmUDYswuWGnlg1/d1t7RbVp+CGrDZchN1Ik24H
EotqkVd5FdVK6MdrQo2xkn6itx2PHljmyby7LtGPLDsPXermNjOg2JtFvqr5IYgfP0TsuLumAVPZ
ZwH+9D4D0EG1hWd4ScEcgpfDamuFrmklp8+OGeA8xiP71HwX67g4jwPFcmIQVmfypSiyUecnfXsQ
xnmOxDYXJB3L0HyLJJfIKF+6tW7WpP5ZH6geiO8V03Pt0Yj+9qFlPtHnwqAGHhuu2kw5SfPTGB2u
b15oKcxG4DG4iccq8hu5OKQfKBhRJQqghksxLqTUgbIgqI36jeEV96xN/uUrgTODWyuEtR8KhoRF
s53+P0tl/Hb/utvWu0DC7W5faoG1NKYb8wAWENdfBwHQehdgoz1Mnf7dt/qFcM78qYBpACi0LAEM
mu4bjG0MEM8WWOQnQoX6umAI7UFoZhsbbX6GuSpYFb6gSktsKeG53jRLvCeUJhX4OeIzuMqpmVtC
9LJqHbY6FGMSiE8Pi/nidNov9zeo8oOEYc58TnacabgS4f37tASuzLF5FTndXPYJS96T2afjfPJk
e09ZesZxbqqUuoLwt/tsFSRr8xK25xh+9vqrQidQ9ldsFJGjxsW2/yM6/LwkZCCVLv+T7mysKU/6
2Y5ej9dw7VJjUZq995xQZdM9GPLI/hC3tEa/jotzDJ32wOmMGUEZcNz7/GoZwplzmR/ZVy1A2tCr
QeW33gUf3tTaE0UjOzKiLuCHBo13wpg+jwYw0YlDgY3Wn43vmxSQ0jnlTxu1qIe7WIx5ihhUD/+M
IIjyT+FD+gMaT9CiRCff0iI2j7dZ6PeJwDEbcwcAo6dwYF0uk1RB56wnbSyA/pUCNWGEKuyL8wTJ
r07aSRZiyVvmNkECgwO04FE0Ge0XGI11Av/2bYW7/wkfOK7Qwr4tJsvKD4KreWUrYothymOwkhHM
cCqRGz8AHc0S2JXPS15Bl3bg64YVJVEJtIzGzS/oyV14B0fmFouHpYxc1pIX6uy/hOojg2kbIhCV
SXGk3jBIUDCLTuZMTIovTVseJ7IREFzAd1zf6Q7QrGMUEUKjnPMsZ5py2QeHP+5vpOh8nXRJHCfs
iHzfpyF//xF8JUeYPGdoFZz6s+DeYDs5UmRFk2jk6J5fVwMv4akcCDiX8uTCBMPqLwZhsYDJ1xZH
zw4Cry63/Acbo23dz7mZbfHIBnFc2uGxt3DHT1Euxb1UrkShbXLY9eGFg+O27CXxYf8PbGrQ7vOK
NZCXc7+URdiSyQ3RE907hXg/ZgYaQb930U9tq+9AnXih1MtRLgXTHFXcta5ttSwToZtdsk38mbUd
zqpsyEMOKNEITUM7CAjpahAvpFWAGDosOxo8/Y+aPw/o25FFRqpGybmYHqmRAWUVZsuWYeUBrdIT
9UgmSC8jeS78vDY5V4LxAEW5xhWcZtuwqPYcHJlwf/9dqEZPQ6wKFor9c/janini/cbNL5ARUghF
6JaPRMHWjtlmLEXIaV2xhTp6qekM0UPZ0VaN/B5JWkJKVkdhlGjISLUF4y8lOIISxsI5ieUf3Bjd
7OCZ7ThoFbBtfThpNKIXFidcrub1pN3r7CXfCTbmKyGfFossgIVVPjTbWs16aAqJhNSUpsLfMIic
kGGQhKF3cNSEjP+81fcAkQORld5YTkoozq8ishwipnwbG7s8QBTI1VZ5YUZyuaN0gqGwx6Y6qaDl
W1dK1teZrxpgW543a6B37WL9mBKwTwn4xHYNUTgkr1mPBlzzb500oLRxRF+wiXavOysUsMlt/GE6
+cUuKkk/uF2ol/uIW3fYOsVIEUdVeUcsHhBsYoYR1uEyUTHs3CKMRH7n3kQq4CmUcOi5P0HikoFB
o9y8Ix6QknelCGMpy2y6AfSnYwgDs8vCvd+Yo1LWpNx3V8ws/VVq+O7lhtESMQfU/EDfYUWyNm8T
8dytoVP4NljaAzk371qMNh3ptbQFrh5SDgROVCcUIgzmgIxuOKH4VjV9uAwXyMkKrQKSNXQrdMWl
qS83o9eIP0CowhMQM4xCuA9KxTayepjl7ZEa2mHHEt3JbdQgPKknKuF7xfFmLjS/Ivm/SE+tyUuS
kBRhR6gBa6GWOvxphugNaWhq9Qf0uZedkSK5ea3jIDHCelSoOGgOQc62HYjl1fPGaMLPTpead8mQ
8X8abgYEhXHDjh7eisX6p/R5uQ3iyVYHZEBKHIYHwMZcZBY34+sSFOD3EaJGrZKb7bkkuTtXISyP
lcT7HB6v3tGkzZxGhZSadvXbQHJaGC6fArkaeqYd7z3Cmu+bIQBC0Q33Zt04tB3/EJ1HiFXJ6OTl
ZVDf/HYiepsoGZIFlo86t8U4iSgghwlfnpurx/JbvfOV8EQS0cNVABKcfi6PPusAwKweOW4M5W1l
heFSKcHvEkUFpBnZg1qOcOwN12pqUq8QavB1VL1n+vz/kPRH7aHkp4ONGImPF0npCF38USsxZNfP
OpjqjsJCPUYX4M5BZCeaZaCTzhQyVvl5GJvaOc3+R3uGaVYR5qdjYqjJaScVZbtsnS6HnMwaBiiA
z/OmgGQtV4DL43H+km8703SXDo8K3X+MI/hZrcR6OCA4quyvqQdaRHUcBc4PafoFZVweoQ3U9JZh
6qMjE5H2FRUIeLauTNu3+gYNdKvy6ftc/qw0NjEwshTMM3czsxYAwt0vroUoz4JpEmbNx3Tnivl1
TYOMxADkHGAl+wl1tFUm1vyYRvp5SMPLizRnp4RSSwN440HLzPEBLe77/JU9d4qBvMzK0o0r/YTc
47IbA8kRe9sqbAmEqloz+X+UJPe5ON0xJKw5COLGdYFmxSvpFv4J28t1rUpC/hwXxzrh+6lFoMZ4
J5hEedl4NOGS0X6SnPRldRlZk8ZRTCGmdHkEXqzO1MGTfaPnLcklTLLDjqvdJHew/DOLkGaxACWe
JBqY9M+4bUHGW6EE37WD9bccZoL/LriDtfhvOUr1+0HOSkdek4S/8YiwLOq2HxOPESVqtJVaSajt
FLvywcEU90hQy1/pVsfkBOFMC1JcBfaO34hL/vETizzZkOaU+HQhyIhJzVZTkX+VGylntNIENEAP
XRFDH76PJFAQPrif1aHIfpJZPjWyMwxssnT2fitP9xy8JtGHHlfsjLIE1lc4ShjV77q2QZG0dzHC
ZeJ/Thwg14EDAXXRt1/4L0WNy3OvTsUHm8KjPQ0cQwo8JksNx/cBHVSLgWkScz4ZNzAKt1kAAB63
/apsotpdKrdEwriwvwrLWJvMAuAbKwqK9I6m1lz7Nsu7h2jpXcNASMD/m8ZKoMsVXTLaRvXE1tOh
KzXAz3ZqRTitxx2gA6LY4JnFIPQQQxBF1dMvaOb46NOQuSEIk/NCZan15JGNMYY9/a3Hh+zroBVR
GycG+b5n/Xrvv6s+jtso4Ct5b8xzltTz1Il1h/u4hTnlubX22hU1oWeXnpFYmMlPlZxjYI4/FVBZ
5hJfHPLW8beC2xXWeDBpjUDxZ46KfBsXNmyGyVqLYK4DCQx19OC7auTA/oCOB8b1TvTWkmdD8WBJ
ctofxl5JiowWmJ6EbQSqPA8c4LoN/tX9i/om5mU5C39qBcepL4R/IelnJhaBWCqUWUyTi2ji8kAM
SFP7oMR/yoelzszU4Q/e2tXgOD8T90+4hWn4m/Gcfi8rZ/Vm3/Wokko3/AqO4bWgWq8y5BWWqs91
1rn2pZQXvdgM3ahqelfpqzIMXlBGKsbxZWg3JE90iQtPJEzh93PD1RK0LC3M/j7r0f52VErCO0wW
Uk3BixGgxdWf7/1HRxbAWqbsUDR+3eYwpnQjFYEpjRmr6EVQaEqCx6OHCpfVhLbJ09LuTiFWkakY
itozB2CO0cb2+HiQUlWT1Gbr9JCEyBSnU5lKENdJ4CHYWerEPQp3zQQkLBI8NW02cs/rEvUiDr1i
6pKrmWjXjEwuehONQNI5CS9tH9X0Zd2UNiMcwaPq0pt6KkkJUk96AJYX1EclfaKfURLxvKfcTIjH
ESCXEKsKMSB0+/6f+foO4LIFJhv3zONqILeaJhaevAvr4PhDlFZAPV6mEyuYDARZQLkBIjuSFiyb
xBKcAugvmtr0rNH7PZ79s5QoRhTchG3Znww7tSVMCCRRIv9Zrq5aXOyqc2XEU5OFOUYooFFLeVJM
KzDgnKo0azT51qIbyzKFH83zzgieoNXObabRy5Amszn8WTxNuNGPNhtIfXVHH6WeltX3HEIBZYUM
HVEJd2zF1BRUUY6Xb5ucmX+0uKgp41hA8Wuhva7qRg91UBqvrIp2oE9bPK/wSwMHrNA9cjYU5fjk
foc12yar4u0gNXpYdih4wy5i0xnA9PGNRibuRXqp+Ktv7oWCK35+PqsUAzTzOpFl5DUPc/Ox8NAC
OuSIyYC+I9WetpSEj2mPgHWZznZDfugU7ABA8zPQBzszxvCqk4FLA2Dmg5fYQ/bxkj8NuUh+gtOs
9DsJtKK9+2b38d5M+FAiRtWc8M97esuX28XS+he+XH3+ZeAKmAU0mglLdZxYLLPferpxBAlZK0F4
piHINJ8hf+1pZGji6XDBogzWyFhjFRvG6nDTB4bNXSWqOGpMipdk29tm4ZE7mbqxAjkuPAGlbmjk
asaoMyDHyN8cs4MqBCkkXFbi5xYxvJP9TuCn/kD+XVTt310zOHbOuy3ifILaSVIAEEgRexG6Udfm
PPgj1YYeVdD5GzPJOIuE52HR2kNQQnTC8IjZyBav1q5jAPKYSElO1UgoZh7zSwx940cfw7d0wmUK
V8ISIlUBGnmIWjtfH8rp8Cdvz5xPhRjfM3djnotOxhAlXnl3SFGBlEmN8ZKKgzyq6J09ZUFiFFcm
pr1q7zm5qfiVZyDZZwDl0EIyDnh+pxkbeb5VEhdcGzuCIAxN4wVAQPK703AhDi8QbQdeLfPGl/KI
XiDXiJKb2IFoCRotL0ddrmL4hNwNy/eIpprp4dHhIwsOQ62f/QenEHTj0YpY8AfF4VIwB+Xtwabo
5L1dyupQa8FgtZeLpzQk2jKu+qrwt2YDSOGtaOSqIKJO++iOAMTumEk2cbAcDoCCeTixNo9bdv2o
Hrzya0YNAIetWQciDpMFh5m6ecqb4u9Gpx9bbgbnrYMNlQniAFQuspuDQ8JQcemgOknmkmlUSqhE
ZPowy1whoNgzbo1QmzseBF64npDfdU13NZpZa71dc7X5xkX6/A1u+svpesjsujOc+/omkCjag+oQ
G4CXa1hEDcIuNg1N0KISONLcqB+Rss8H8MPZ5vlUVxryOZiyWfmx6ftq+yIPi6vXCLXZQzqr3hvL
WNQB+BmcA4ozOEEruG57JXP/b/frYxvlmFsxEg8fkwlfETwtpd2+7hBTOtTwyMVtCg8auN7plBku
D+fwkVOreuA0aUHuulyi8va5rWe1yvi8PvdtP2wMsiJYpEeoR5ICd0UnbbUJGC/J/DS1wgYd0Sm6
Qx/BqJoyudoHIXM49pO0tNSbNe+nv83w2Mr1VkrvwOUvnoL3TLpRSMAMfbMNHhofC8eFvWsgmIxb
/uENRDyXzz/A65iA7rqMeGzKmm+qso8tiw+aMVyuUIhG7RQUIhhyhMN9e8djLBhrHXP9uLz/4nKe
lZQ6PkdM9LWXg1CiTr8GDcLumHiKpXSOaCfM88hm6h8veaotRz1Y7Ko0xbz9qNaBC8VwCFp3KvCQ
Hw7YndSABy967QBUk8sQhSHKWSSC93C5XaZmu3Xabfv4wl0YMu/UGZ5RWVhpT2KuwAMXcVVt5OOv
ik5n1ymy/mYitE1ip3IoeireLIDFoqkouB/Bh+m1mgvnWajRJv/0E/cpG67sasQLkm5YJ089l02j
LgEJASeCaiMPPHCPD5wF/3S4q0SvYxf79XhEaEqhzMDcD5AtP1xL1qVPO6PUHOp8LFa5viwZLTtA
NMpRVYm8G0XNyd0C0NXfdm/gfZo+O/bR4AbrGD7fzA5w8I3+vphv43CY4Cw396AYsYVQnn5MxdO1
dqDtCpk6HRAheGGlPz6PemyJmxSQtNT+xRVfOY542imEkNgqrhfBLwlP7fDB276eaGSPaoftxSnf
wKAajuVAoiKCsgKxzseV2n/wPLuulPe6mi7hM18tpSFjnO01cAvPev2B4XdS2jwMMssO+ts3qv0G
RS8oPnh9+RnICkBeHeBTABahG3Q0FsWQbRlZCJlCeVXDmhpjc8oXUwbT2OtfFE/o0u5Zyj+LT0T5
OhA9hSoSIo1t0htJUsx9erens8q8hn2dgBvlZZM0gDkY0DDg86E5axWweQsi8eNvokNT50ku5DYk
SKUI8ZTGUBlh866GpmIx4jGDNFsZNgqtNNjC2yJdrkupcCYXQxFeCla1DjSFDpxnxw1eqo74KDoD
M5FTxKeALNMyvjrw/NQpmfDKcrG4dO98aXotEHJgRhCFRdqy18+C3poIO9rUXoESLUAeWnhqc4YY
PZTQRe7XctsYs7CAKGUZDVTfRe4EyyEv3AusP3ydqr22JsGphdxRXxd/g5dd0j+r6I4h5k4Eu5KT
vIJr6fZTSsNMg7turUm+e3/n2nf2FcQUDeLrOubd5x6S6ZdYHxQWooLzNBJ4BY4wpnrJNtfSIgxa
XWbVYCbOc6VaC8z5kVK3ULQOUmL1n80BGpgRsd/CWfoHUU8w/4AZPB4J324IZ5+V9/KdviV6S2xM
j1pRF9ONPLqsJQUWlpUmUIS0ojI9GVaaMTm87eVWvRVXf+Pc4l6tmryai3t2e9uigi8l4e1sGJ6d
qCGhe4L2iH1bApbydi+ySgeEr5Y7zt5H5Spn2ex1yanRgPaB3cVxr/G1PLzpOw2VunlmB0r/jqUe
lPe60JPwcTaAyLJuqRYVQu/LOvLndA76u9bDWUNHxcvVl5L0jiVrv1uBZSCNdax2hL4PoEbZsJM9
hsxnHlDMs6z3NLoKgWwWwjaRoczNqWC5p+khD6n5E/5x476N4cCCdLiGuyzXpkusbrck0CU9GQiu
+8lpAbL7PDji5JzLg6ia5BCKyBVy358+Z5eviJ82oc37rLTE3xF6m8h8ItnmgLmFl/6CwGJSL6Tz
R+lWCgsLgQkrVD3t4uALuUsQX/005WoiXixF8PNYAcDCLyRe6476fb5Br3bn8aCzAjIic/hDHjJL
vK8AXwbhhHZJKhE3crJYJ0ZK1S4ipXk3pFBIWfaDOztgA8zRU7CIPfasFSd41K0HuQYEqchKX48w
G8y8QfRs4tKvmhGFX3fErXK51pTGNk/4yp8qg5qj0Hk6o4WtL/79VwHry6B0m4qjjO0P+zTnK3ck
L3JEeuVZt6czqbreCfIzW884LjaR3wiFL/CO4u+83t/zxUdhCBGq4FbHr2CSp+3MiRdnqkSofyi6
sArBpPCjOBVZ8tsJ3iSz0d++46T6uKK5XEmc8OnjF2ZFwSC3nCWfag9oq3xP2bJ3JGmz41lWIPgh
qp9uEbpADuzEwhd2uAgIpA9NVat4vOBgcqcNP+fPj4rLQs43r70twVLggDdMHPDFoAivJOIjz/bX
QNGcdf2cLWFXz/KPxY6CKcoW5rQEDUREJ9UL6vIzMnkySmPwI0pUFcpHYaB1SDJTb89ihmWEooeQ
evrlA6mZ3lmxb/keF79KCrdaKQWHKF/RTFYLONvsqX98llSJSwWEPKiyAi4Ub/3Mcwg0J+4XBlwC
QMvAZLG8mo/Fw7Nwo0LLTTFI/vrVrbrhB1Qsh8EKi7AvZgMQKQC3iO+NraIkC5n08rq4D+Asp6S/
lmt2h2bkpze8CtOVo7IUaCo0jcGaUziop9YyD2tI1wOnEy1bVTXskwJ6ygMdtD+1UkCenzAv+yeK
IQmKQr9CWjYtv7u8Gr7XtUBWT6JsUiHUvQ2DEqmYHgo2ZMDWKehYoInSMeZLIsfv/1P5+7kfDwTe
J4YcTnAP5njHW3+IcXraurmtzXwn8CKv2rXKBRAjoyimjYUxbAZ3UxCl9nBq+7VktOxALvw7YrNA
dLLXop+5r9dbRd07xq08hseYsHqYOBT/22j8Nui/rW3hNJsOhYAGjjT3btKIkBpT8LktXpsopJVw
nT7RrhvkE3hw7gpQ1n3FcDgAELx13bvNMykD/ApWOPy4Hjt5aRQhJSf/76u3wcOnUek0njo+wM14
QBUExQCBB1cuD6y8sSqHbefayqnb9JJSG+Vnk8Rx7pOPTkbghe/Rc04EYAvLyd9lnLguUBYLDF1V
WQZW4jqYZ9vRApTARZwvez72rgQIEP9NlcNdO0xqKPXylwNzDmMIN+SpptGqx3VW8cPvi9DAXZFY
iNvc7njuSyBNzKDMXn9bDnNTZQiEYtBUFPhsKFpiXqwonnHbfEx2sXAtH7qxZxi/kVj5Qm4ipUeS
xXM6NkZClYII6fsbpe0ohkINcs4qsdWaS6JTaaNKE0tvNe4h5+TjNtZ6oXNfcGRYcPELJD5gdTFu
KqPMTTr8q7M48xi7PXoIA17Eigiqh7rD+Xl4CO17vpzHEkVHNBCStG0qhtZH7UiCDNLXPPriR5lp
cpNmf0eth1B7XImYDHAT8lelx7vn5HdBmsf7gZPojEYPPLbfZLF+Q1Nd67UVbeGoK19x+qsqd9OI
x50y4XCBpvwBL4xy9m96PPBsp5exLXEThn9oaEmul1SeYQQBw/lUldjvnJKj80S8atXR9IFbodow
HqB5jtE8rW0Y1TShqg4wc0Nro5QWwwNPVuVC6DkHEWnEGHu0JmANDNXIw8bodFHRDXcDM7IDzV1o
T/uxCA3Zi2/WMhkmqbkq8rXoMpM+RPMsuhNAWH4cfwOldDphxtCZvJzW6OF2he+EE1bqyA9ALIEe
6RhxCIXeDjZoUyP3de+1qDQApfiqizpHWRBQA30+nHKep9wfv+zmThhzvusBoXjuCLua79wUVmlC
vYytq7mrStrQeshiLv84lagrXa6sHfJzS2hWyJw1SlF5QZS0hE/rdtjqK4q6s+LWwPVh8EM1k/sQ
RHmRkSHqqf94Zi2ggPNxXxXmED4UNrKqgz4LBjW4LPESEzWqgXxN4q159+YglK6F5NYmmDqqsndJ
OQ3azvz1n0056fS5Rk6eLSo6fTMqNd9ApBqhBkCM0fRCExG7Z2BIXodh7RC74SjKpxEQvwrb4ziG
kYltM3xZasaRh81/4G9VvJG4uWau8Ul1ziNNtmhPOhROxMbW001CRB+bfySm9knhI7EhCoPyiAk+
Rm2U2Dt8m83VgWnXwowFcfqCwvCdfWFF4Dq1jzOkpYshgTz8HCM/o9m0xaBfI7KFkeNk0UEDI5+e
0OdVyajtT0lKm/7FAD5bRBtLxnqoQNSyaK4Uz31sWOwgeGHBSNoauzIixHHJV5ZuqxKTbyG9nWJ2
4Twf9JFRWmlU98+1ak4UUQzeBm9iN/78hlnRJfTPeV5Umlr3YWqjkEsevfKqJBejhh2L7yPLQnK2
HLWshoQlnMz2zuQnEfkwz5H+T3L/e8CWqaOg6Ex2FMs1sjtT+DlJny2gG6ONa+2medxTc0LGJh8k
0qQwoGkXODJjfgX1dtGHuIXuv/mbTSbkmSF47bPxNEJ1nzQP7rZeSTG4XOE0ovogQ+OhiLpHxnLq
E5IZgMcsvGqv/LBo0W7tXJ5QBqeumNLkNWiiRTbZvCZV4VNJPDl8Lt/MzVuGoZhTJR+WGqG43q+k
w1LfjnFAc2kcg0B1y2Bzv3PvAC5pePrXFnNZ7Ht77Pt8hnfh/Icj3iTxtd3AlMxpFA38D1+gDrib
peRZmqmsJD+m7oCOvlyDflmQdLXSSXo0w9cct8HT+oH89ftA4tMsXqIq/ZQJgCWTKZQa65JkpHML
rgxiyYdnQ72i87mSVPIZDyJKIVTTgYuyW2M1C2qExBNpmNfOYe0laSnQM6jrqPkUEnUqxC8NNl3i
QaitvNmkR3z4tUWdpc5qzLjlHStXBw1wtL8HW2LDXF3taRny+knMlIY7iz08FIW3uWmSprKEdoyY
Pq1h58MYm6FuFyxb7v22mL8r2/4mKj92wNXvc44xy0lM0z7txJuwm6NHm3/vDQOTS7vhrpVxb07l
iK2eKqO150rMLSUBRueLjXFXfEGq0IzIBV6/EIO9840CiSCWY2PsQTijeAymGkWF2lv3oRgQtf1b
dEyR6/9m1kns/kgPp3K4PYtqE5j7HZA7eGvmoahwBQERIUBiRRT9WpXnU6PaZ/Yw0RX6bhYYcZec
YQpgXB2g2MwRETBvYYHDfSzg1IggJZjMTABU6O4ZcSHCALIT4lwMRelhtLXgdLViTgiv7NgyBkeA
lv8ktxd8Rqb9xelfCvYWui9FOfVUMUNXa8p/K2ax+48rbhAg9cARKygBFqgWMs12r/t0pBn5fCLY
WLNNoN5H1QfR86rheG+p4RlA8IQdw5BUge/pptT8seN2mSRMjxCeD7Gy9Vef63GJskci6zn26ESF
cit8rKUpuL6KY9Y/pAKOSVyAGPKy4oGhlZFIYro7KnYUWlzh9JebJMQLFdZ6+vbutixo0ukeDplx
YzWMatRV2+O8npb940qvFTZWT+SO4RR57t7DaQPJMgQ1MgfWTdP9It3eneZ1jiEuTt3Xvj/i0Eds
fDz1mWbtcg5gOGginsZYr8+lq0GeNVszwxFO3r3CSRj7uaMuZpUAGW2tHqSP1YWJ65vSnPvxu+rQ
nFxfe1lYoj9JZPnyeSmkWiJoWi4OqiN5gblARPgjue3i/1kqnzmH6+9TMmhjnvyd4dWT4wEfD1+T
VfNQefQqOnpT/oc7qHD941kPKO7nfHP6RX1vrJZkEbjTPZE9KZlZRWM/M6CCW40lqp/rDd3scRVG
5WTpF72gOF6FhdswfLVHx31gwFHLgKQ1ANzQXPW0Ujqa6mth7LfSTDuuREbh6G31XfbXBs5REuPW
vZxkKJ/VY7l9uMIM0+sHhqjhNFuEP5N8W+pQNurGPuOp5UL/xfnCRZndawQv/AtuiKqzKEhforw/
jtrBZ0nfaMr9ZCfiQwr/ApSzeOuiKFcr4ipgWBlpMgJBqPoVJQ11VE1BpnSSKXeYRSsIgCRYpIRY
hqfXFnISx62DcKF0KBYgQNDIP8m0WiwDB9gGMB7TU7r4dVuNJRqGdhVOLQJB6ceP6vj34vdTEsih
IryHmpeOx1d3n5i/uQ5K78EtDvSL+uZrWO3C0wNCbP53tF2n72uJZBCaOhJ6M+Wj9MM9xku9yjvv
dzYIwRUFduQoMn35DOKivLD3KgK9aWRRdAxrEphjMePB8IFIThtKmQEIBRes1FvZ/s7hckSFGVYV
tqDhIHhTOwwObeWuJ4ZGp7AN5S4lh/WpcOsDw4T13MCz2ByF/aEUvLXPM+KrzJBQbQOOuI6ySe1u
ujPNT19JppunAK20L7eJgQMxuxM3AqO93k9FME56rVWZ7M7NNtWrLI1fyhW7YFckBC+eV7Bo8qkH
hW/MwRG9geALoEzYujHboLf0gVbHU5F+bx1DIMOeEZeRC5jQ6rc96vTfwseYj5ZAD586ys30KQ0B
e+iWQbmFg/Ih0B4Xq/K4Pe3B3Ln+VZ0X0aFGNyhs0bRpAuIVOjThITiryo9v09rxZYONtaBjHiOx
7o/2m9+1V4UG8pZQjK31zBxWjnAj2/xZS/rAOSDBsYzz/nSNswfM15EwrU3Dp+YF/BRTnTxsJ8yT
/ZJGPGc4vezK8hQ8AVLjsAyJsrW+wfvBskNtMPTOJKZSnPi1IVPCpIBaBO7jb/GfXiD3YLBEo1w7
aBnm51qHB3Mc4Ic9NCBlfUuUU/G87OHshZOydnA4pg5A0/BlY8uzWXt0Tl6HscvUVUKGsibQOToS
0/ni9KKogYJD0klSQxT9botk86VmheGxsKmYaQHh/z9q5VRTwQdRPqnzruFBBwgxQ7oMNEjEJzAa
isz86M7gADQNyEtEbCTKQeBY5AVAYCek4KCr+c9aQSKxoJ+pdg8kx2bh/dGTjROIiaApON1wOmAV
8aBRD2DvMp6ryPOEJ1QlkBxMpzvmFf9KxiG9WOlPbf4yOQNJ7lQLvCeqltCdGxSEgjk4qHkhTLVw
5QBOWnHm5P8XO0pe1QDNvTvFKpIiErUS1v8rKuWZMn3U4W/dvc2rl4DBustEa8sMVoJEy5BokrMK
emVemEefJP4qGSPcibv2u+w3nPBRVWp3Ysfk5bM8e0BfjlB349XwezAdRBz2xprLCLOiogFCKOY+
VqCRgoaySRx93Fzth7Jo0HGOFNQYeNCuX6w+H9GlFfpsBcgtU1CjDthHjQPTIe4g72Y5lgPLoJZH
uoN5n9gK5bn/sOrR8JnjqAzeqeCH7/3xTDYGxPSA3idijrQlt0jrDddsmGWh1prEQeyq/Gwswvhi
zSRWXcW4jb5KfYkakC3flbFkZ+0XVkgfoRM9TU5AGz16iMrk0W8t8Ij0SJV1aIt4LMAJCbbdjEtC
YUmCkmeTzfvbXSumgYPaNGGl0MTsj6WwH7acbqKaNcPlv3XMMKP4KX7CqvhsFCforSRxrnFwEgQy
+KSUh7s4PNWuZqyUh0mFMF6Hl91apdsr7SqIRuAHJJLQG8kVw1zwCELeoFPwnZP4gkCm9sq0k81s
ZxsbrpMslyzcb9KvCDyhndn8JVm0UTFjmDUwSJoQBBxZX9JD/SpCIm5YdfYZDUT/BvPFMRq6xGmo
IqaadbJic+IWJVVOwzoe86gfgBwun4LYkRztXmbcji0sYaV4u0lcehauRWoAJtBw42KpBvWc/9G8
csYT8DGdBaCxyU9Mje0fY7ho3MdT3yy9t+aVxyq4j9UoDfaXIq1PS/+Y7br/Ju233QPlS+VVJxRD
HUtaGluQIXi0+A+Zk3K8eKI6kKm3nPRp7En1ELzlWbkwvc88jwx1yRKg7OFr3AHP6elMH8nUlkwd
spk/s4Sc80TNDsmb3jmNHu3LMMrr2f1pYZwCp9TGBEzueuHQR0/vEbqVkqfzV/sKSepLRZf9guPB
jtOs1grZEu+WzZU+gGorQ7SyLHPj8bDASY0Qmg+aGYAA0wG3jiFz4BmveIHw8BWDerWIO/c7c628
CEF52k84j198XebOSBNjRsNy1Ad0L3mqQP1bRlJGsmr9VVFYVCbk+pRl7tfPjb5syF53uJWvWcuf
o/BLuAGwjoWckwDL7dikRDSEv7Tk0QbP48mDXT/N33gX8gqj4gnuHcnc8hf0PN2FpxDExYFF51XL
MxIZgBxCDxLncKjudfiOXrl6kNJK2pkkJuYNor6suZOKqu8VdNo9Ug0FBahG3xmfIaPr9j3xUwiy
S3ulsdKRKRtuo1dJOFulA3ttQw/Vp44FiaW9BsJx/Wv/pBMH+e3AZye0EmeKSPd6PFlKEyphIF9p
2x7PFd5hEZMxjREjAo6qpHjWd487iDS6H2b56WG4vAEzLnVoB/pIERtM/eHc6ggI/TYaPaBrj6PM
sH2RnCDPs7T+xR9PHs2ojBIdEDDG5zful5N/xeFp3/dqCNsh0aYMW7SwvMHB6UG1t8bs+c1o4Muf
Gf1fE0D1184EF7SwNsMAaJxzMmD29F0cueZsuK5Tfqpy3H5HgKyitnj++1lAdqyoP4z27bcUtl2c
a3ZJAtukxeNpXG6uLY6WP/W6Y2ZRUiCyN5FY0+O0qBy0jqzBPAHxL2p42mMSjPQABOWyBGbv2oBD
ZO2FNqyKUs3wigIp84iOmzDaQPOxPHzblwtCssmhCpoRtqxIPAv0TbUhhRQFbXqNoglIze4TQKMW
D/n5e83Z2pDXscBLdKvIifAiuvHtFmBF11anVat9Lr9YRpPqyFqBkkAB5GQDXc9wpDsitzXUj2LM
DhcG0B1QUzfmA5WwGUwk0g3gL3xQYq+hLRdv1U657A/jJtVc/Y/iE5k4L0Pn34NbTK+DtAUMu0BI
EcyBpkS7uLHoGMeYeHSjToCXWnw2Rx3/PDsXRW2YooEYBKnzmD9rVAPEFFX9JYsd5XwV7JpUgFUU
bazLTCh5lG53fhhH176iJ7CoZabVeUY6GyJCxRwSvorSmwp8BBDfz6tJhBo67ZXQ+kJFF9NgVw/h
caxfr4h//3iAu0SHlF2qxq5Sk+f3LpHFTvpXF3SC6erKVqn3JM+APdO6oS4+UXnN1Ikmwa6uAcqq
sDXHxHVUZ33BZFBE+UGoaPRDbV5pNJ3yZedW/CA9TAB85Q+zugaFJDv9dfurixEycLTtz2Yt+9j8
xuRgnOZLUVc1Iiv+PXlp0bvAPiGEsg5Iryec1mOIho5WSOky/5Xe74vhb/P2/brQQbEphjletijE
k+MjqmNJmU4toOjPlofo2ToHWWBmtTtUJkblYBHJq/tnjCnerNi7zx7Zbg8JcBxwGnu+O7tdIehT
mzSUppl/z0nkVPnR/LQud7FSQNM8FE5EH8XWQDfBzJRnBcasRhxOz3PcNUz6hLXfThrlMtoCbdER
w9LD4fBMR8sEwQDdEgx2YANh2D+IObfptEwV+l8GIXhkOd8PVB+dlWzqm3La5ViAt9+g7q31YQeA
4tr9CHcvFtwAjet+RG8Wixl6sn7QukRR3rjRiH6NxtOoey7kCq/EsTUwa9zaJTVO67mK8siFXaPE
ZE+UoLkSyRQmPwlFoDvVdHtmPBRVIGUzOc3v3pCWYZB9+vWZ9/79srySu5+MjGGl0brXDdPe6PhH
X3Ukcc8kqQdJJKUk61BKMng4bzvdfcZB/YByKG5zZLZdrmcAuu9G2UsDVL8qj6/zjdc23K49oUPe
RfcNv1buJLIkpvD8pIiPGXaJjuFsYY05OdLRFHmdA7N2K6hme3ljukv7tLkiozQXuxkwbCiNdu+2
iGP6z4iSrK7IMQpEgAI1g6uZAtM8gGE21ZY3y3sUneHDsmOx+oisd3qJjrUTiRUy5UyUgCRxAuHr
2Xo9QqVq6mwH1mhkz+HFuKIbrTqUteyIoPZ+u6e1xoH23s5skq4vqb0p7KPUJ4DQ286G/V1Jr3EM
bAza1IphyXcMIu/H1S16pFgGeikIFeafXlsVaP8QF4LKtcWRLzDeyOxFLMkfIiD9L7P5dnnQU4ST
q4EhR1lljvIoHiat9gqgdABuYEuyDYZykVLkPBBT85dVj+4UDBbT3OTwC1im8rRuG03fmfc1+kxv
UGiU5qtYTognJtijIHyWhW4voRf4MBtwg8J3WWF2a8bGX2EPB7J98GPFjIa0D6hSOHHzT/j1uDoO
J9rlf9AzbCoOeBAO3R73nMqTP1RYriZNELHVpaaALOYrwFfI2NuNsP0Jc4NMfrpN9192lOrirOiS
6wIgi3ck4MGxZ6i392r1oW8Io/ZNrGrSk+pT+af28+bqY6uz/65oKnTjvpXFxFHQ6p0ZgA7rmfuj
eeWpaPNlByCdvzObNZtfwlxjhXMo8C80h1XGA01ZlAaN8E+AuOm9QKXoG09DWHDNA2nzknz2MA0N
s1EqVsV/Zwx1krKLQ4yBXSmIHutInqCSPeDytb1THifvf8lyg4V6rS+sg/fI4BcjBWv8F1SnR3O1
lm2ojnBXpmUfoTwuDPoG4U0kkyG8LbUU+AwtweOuuVrmS+4O7tsy7XU6j/HEVT55SbQvawbRzd6S
kjeoWtk1uypuSjBxx5vngKgv4XSGkVwoF3t9nU5ptZHlTKhyxFvbnt2RyZcIvDBNmA5OyR0vOy34
IWjPnyCTE2iRe/WDmmIQP5De+Y3fGgIXn2cwqeci8mIoGrsoBAQGny7lHDj5TFOQn+Z741siUZt1
rB1K2gfFDOgfK8Y56eKxE6kb6CbqnstW4S++qy3UYVjhLyucgij1feHvv3tQeS+21+4XCFBXlGY0
c8QNg9QxginZcO5QbvN6D82h5Tl0GoyP7mPXep4Mkizz35ExewxlFePFOCVNtGjtsm8sexEOayJp
pSq1YVpdcHm+OFf4RinHFyEV7UNp5JYZARzcrWEU2yu/dPJ6M/6kwy0osTJl/3LfLD/77dfOz1a3
MVMEekFrezOAm0guybdB7nIULN/zJI7eag0EuXLvARcd11/clfs80SiLw+06SMTNpdV3aE+LqDMs
26o1H1MN4t3ZuOqcTCitxQKnX1Rz5Z1Sa4zSCayi5YSRVqRnix4EoiwRUvrBQ+NE40cWBmyZ9NLj
odvJkLdaf6HAEpS9MZM3jPZCQqlIYePVTssVBWO01z7Y5gUD1jwiWV1X6/mgm5hJVdT/lWzrh5hK
Bvhya08GUNdX+OFErBkJ00+pEO6XsjD3A/Z4PP00wd+7JDQ/GAZvnSs4y5F0AzRa1HyG7QsY/XsR
FlPbvHMp0jOb+ZZgIos9TUDyVc6+FavJwgKlaT7zbHamR9LfURiVQDKc2AuxHg3pSP+SWCAzMSKa
DGFefA7znP0gYgIXWjjhTJhg/9ESV/Gi70R3I3PrjbIkO1nbYgQf9hMZXMux80rZtMBwuUklp+wg
Yf8nMTA3X74LY1gQE2NlhFAXpufrD+y2zk/9mzGoi1U33SdPxWowQAfmBXDmvAvFdUcgykGz2djP
DupVaXfyzCu6ObGCcEyuoL8CLQQJWeQ4sKsSbmUvtuAZsOObZSiZm8ZI4Q5s+di8Gj5nGnfZptOf
jua/FtGLmtyla5euDSd+hLvt/zAGc5xl679TKmf3HF0uFfyBbGqq5PcTMxmwl91Ls/c0vGjbr4/A
wtyyyL+R0m/OVznxMNFFu8tFoC/T67/XrpJoTwvKIs+T7S2XXCwSwqNL4ogI+qb50OgsVwVkrRyV
9MeBGwA6wlmQVPflKukANI6KWovMlFQQ32bIJz+0BoPYt4+sReX9+csCjThULmXGYXbDzqK/Wsuy
vUGDlBU9/LWVj9EE6Bi/3i8KKeV+uwLt+WnPd6WvQGYJuXQ7K1SxSIqnh1TwGBrxB/DnXMmPDQiR
/EM+Xw04RgZwm8N0BPAK6ETMpfahJ8AAFMDRFXVXBWqigwbSR7eU6A7u+Nc5Wnz/y/vmTkFJLseP
EKgMw39UlIslRicZkPVoaVAj+ANQY/76BG/ohorELFw/wPrJCAHKV6h1DEfD/MuuGJxh9JQ095oS
SFzqKgkcXteA/8iUhHTwTWe7QYOej6ZpNxdpcAodcfaIGy2BGPb+ctbzG2X+DsPD2q3x98g5Ln4S
0fKqGKKrqWb/o6BfKzVtkKz181CZXCqeTyIp9AKKUg8pUqAeeSrNrPRoa9YwzCrM49i6VA6w4jbc
cYipfvnXj/1s42Zv1ETiJUoTRrFCF5vF9Ypm4JkqFjTKiJtLb/zGFWiBQ7Dl2yxMxGtGIjJJVnfM
qFniggGO+d9p25DavWStNEHks8E1AO2sQ1v8d/D883/kdRiodRBARcSYCzFeIkWPewSgUhDwVHAj
9ipJQYpmFEXVQ6buS5dsf9yOYkt8g4rFmCjzRVn+ZDBscpnAxa/3SjD3PvmWEkaEnCytF5eduNx4
2TGm1wGUlcocPjMBl+bohNbudzSRfdjuez91MGrfL2EDZ2s9tPINY0mecgiHG4U7y3LjpARJWb83
GME0ypekMvasJ2mbl52Pn9XhvS8553gWC4McLqFeMaMuHM5XjBrQX58+TBtmK53Wp7wPsNyORQul
lVz1UoncJE4myo2d2OKqWIIJfIH4hBgB/i+mX2GCkQawLx+UgkIZGipfSXkE1jyt88dHfaCVmgTO
cvywTQW6G8pvJoeMf/W/cHsD2bzGB7ehKdFPY/FowLzpTqJ1ZiylyHaLYIaXwFv5IOp8+UFZ8iRs
SjiPyW6iEbtsr8QKBRIZZGKQK9BILmlIQMlh+yFcsOS+3BQYjqK4NZEDlmvbjvTvgc5ldKB9xJwZ
QRn8FCgj38jUa6p+s93dxCj88EI0sOvm6Y8oDiH33EAD3Evjq+wfy7QNQmL5q2negRng1Z9YLH69
TTH6ie6BIpQPFexn9pnWHGPBDliboJ3+O+DpF0FMSlQDfPOtZLeddw/+Te7D9A8GHB4uQZUJN84m
9rt717pQC/zHDgFB/vSPHLsXzh6WUg7Ba6XtDlltmiEHE2cJKvJobdkgOL0k/Vxvfo2aFWKtSlUT
tvocL5/MLtWXMFPebgaWxmQyTi3s0FLFwBQY6gaD+M5Cndj6U+a7W3omULX8hM1dCg0e9QYmIg39
8mpmeES6FBOxnHTqeWEbSvcYQktSDzHSm6JYZXDqI6F1K9nNxedIOuUt4AbRHBYmmjJJKiqMpxN6
InN+z0MQDiWyTxmoWlSbVJwOMoRfC5SKW21hmTGyLODReZMm9CDB8B/2+HO7MRmNf2HH8V4HvkF6
5cIZxVE6lgGFn21Ub7ODH5bqcMiC0TnAmAqa2QTR2HrOSHHfdsTo1P4QB1vOcCqME2jcIMj14uJg
7kVJqi+7RpFIRmXmz7Nk7qsKm7wem0J82FBMm1k5Yv2kZ++ANLSiTeF5r1UzVb3DOOnJRRdsdvD7
KvrEdgXoXkDj43A1ld5SqBAwFaNr5SKg8S8Bono4dPzPuvDZJZLFRdjujUwjGOYJoI/4Ld2FFrcl
D24S/FsTYeK3IM5h1ChBkXuruzdHeJYQIJ6xJyhCJ6aQVKGokapUsZTOnr5zJDuhpS3ifNn3Ckpw
1BWUmSYaOLuE2sbniuCwPW+VOkFMeE8zgYApOZb2a1wfn0yAdq3Pdft2CbyDOBYYXXwI6I6zCbG4
AwHdNftFDvDRApiSEnbJDed5zv6mPwmWnoS3XvLCX4bAmaJLk3C4CFIgdCGj87pty9gaFnaeO+hK
8wuizERtHU2ACaqNnzLFRAkLMqgitZ+DZZq2jTmGt8dYf5xbXMMeH/5Kgyv9Ycm5HiD0+sAoYsiR
j9Kr+K1Vi57rzypZFf2SoU+toiCiU5XBiKRJ/eTm6EbLzzZFG/7ykcfx6XPElBJ5Zc8dZB7YQW0Y
/W493DiKSVRkdwp2cdSK1rXqxXx+MS9WFifUKU+7byE+VD1Qr4qz5e2ilFl9DT4Zjw96pC44DoXe
WUBBKLG3EslmF+U669aT4WWUSa38q9IN87dFmuCY0aL0PaCZhKNf1criLm76Q6jCZaClITUoVBRw
ro+dBQoYtZCJ1fBPiIGZ5sPp5xoMkcUITIHfBrp0e2nhg3Bge0IMkKcJsQOqDobhpDnm5NN3pBFN
zQKKHc7IYuTcGzvmMn6PurCy/opU8YKy7gvRqDXux6/wswhMppaZ4ULuWPw7TQ9EFQMgly6RnSgT
FDno3Fb5DMDN+z9uy6Dp1rWWnuwx/+3BR6aNJY9tbC7gG7b9QdgRFqnw6oiZjAxPYY7fKXMj/c5H
pWj1pltZBlXAz6X5KnauH1hVVGIYHuxNtx323a1+Ld/2UbqEuwwEtcaH7I7I0RL0VllUQEXl1StF
bqrsl3Sv1cdES1ybCScChz45JRQLk3RjZTRO2Z4BbZGsFWT9CpI9YYJIniaxACAdPCnnRdtWQ4Da
fzs7ObVjHX1pQe6IYQP5ByJBxigfAnRiQezZUAzzZSUiISCCKdmCbpw+gN11Svxft1wgC+2bhOSE
CPO9jXcaTSHGWayESlNTBkFS2TJ6s5pHQO8ur6e0JuHuM1I8ZOgZ11IyFMl4dawJrfv476KZoqNJ
gmCowl64fwUEYAkAhMsj4eaAly4A8lmoiAsdm73KuQkidZMFOtz8lleSgp7j0L0kXVkNmPy5Z22M
4RDKEuJr2jFHgAOOFOUkht0IWrxGp7Prjeh8jY74VDsNm8F0P14W7aXOygz3DVtZQHD84ZGixMp1
THyYx4beMhCLcpHX3npIlbcOhgQxFwS1JioD8OnfSYiwUaUxjP9g7PIKoTO3Vp/jGI/xYEzvDyfD
k93UklDaJGr8PykOsMUODo/U7FiZi5rss2dAQfV+fqB+zUL4XWltaeQGGIFQR16MfSjgRlvcKSfN
K9qPB3qP40915Goq92AnB4UoNnBT7WO+hoXqA98AQ4rQaRGB2a1zHr3WyuW97WBUJKFLz1Qh9Rm2
qX+DQR/7C3eNwt6ZraocIphK/yYufwW1poiyI0wAyyq1YRT6Y1DqatBKP3aBprCSU4wGXNrkvDes
KecOr3JrhcVtZRnUBDi90BmxOF8nPSYknzz8+ZiT2QhhqYBfx5+5MFIltz0c09kc+jgGpplsDloY
jfPogY6GkTtnZeoHXrWuBBsNuPzD4omfSVwRhgrW5ALbKAm4eUZITiPwgN4ueWZzeZNJGjaBjW6+
w1319e27J0Nsppm3SLKQuRZNgajfe57+YGpcsgb/r+mTR1RY2HASLhMzY3rMFicKIqQA1c2VBu1l
r0DilnvOQiS15SjZ6ahrk2ADIFZUqsqUzUJPXCLPzEUQoOJ+maiiVUv+4C2p1zbcT0/KYehI1GSJ
amvAgiTh3N0yiKn5kkbl9naGufRZKyV0ODSDHh0m2lHN2AlU3LEMP8IHAPA9B/5HaLdXvVr6Ksx3
mRobPJQjg8z1c3OQdMbZiTWaBHdr1GxbuXMT7QqCUM5tX5XndQZdUMgMkG/KtF6twBjKm4eXHtbO
4TzFbVpG9T46i0f7GhXlgYjWL7kvKJBG57gVQ9wavh1/pwQilEY7/wq8fLDezn7MgOaZjBfkXgL0
ODDxN5SNVLTpkCsOWxEyHRt2Y0NOL3j1p9nhf6THEsmNnlb8p74rYMMbJGrq9SIdzO2lpqyI/tJ0
u/7H9aCNO4odSgSxnMIvqKjMSPrGiUDsuYL81wONIb1Pb8JY4416c7igF9RG5L2t7mP6EioAUa7p
kqmoImC6gCS3K1U5QsQtyc/HFaUgsXHn7qBnACVhoR+kjmbp777vfvWiB2Qc9YMNKZDSfIRTDZNf
7AstxjfZRpOlQqB9I7iqMqdXjfYzbNAnnmDrXgqgogZt7GvzTrE89hQTrDM7Q015DIPM0fUfRDmv
VkAecPmXT6NJ+QTOi+UQboLorxRlaLQEFF5z/rCd28uyNG4orGvaWA+hV2VSLhSotemHIs09NTbI
rZoIhmDUEpWmWTt0ScQ9wdfqN8sWTrBrG+h+aZ2SSapHsWscnhk0Lc/HwrxrWBR5K/ZejjqNvHOm
C2YfiWGyl/9rH2oQGpwe+o2HjgJpVTWnRt222QLGna8uqo0+I0ZFW/Ja/2jWEOJZohCrIvbcpFpA
sCyPWWDsEA7TFu+1aY4TshuyTot8rD17GdDLcmDAtSXB1Y5wcBlXuZWubI0QwBJVcTF+I+ulOlSc
326OGd9+CZ/3fB3Yh0lx/8wIi553yKdct+LePgmrucN8xzR0vO6AHnfIJ3qRKMKby4GwfqoJuMhc
OyLmWkqAI8W9v6CiSls2Vg/732IytIVQ+5LmbJH6iPoc3B59p5qY6Rjljv6VsT012neJv/IPOJeM
IuzipZvPELM6g64fwnlw7B1qhnvEGb3LR+RgftJ7oAnbu2dkoC0+ON7OKPWLHa954yWJTsYI8lLm
9BF95pre4qTzJQQOTWvnAeb/oN/KlscYVK1Hb86cxRDUirFshJ2WtDJVKHl8kotV8lwHdJG69Gk6
DoPKUOr06LdDh2/ddydy0ypN89DvuB6kgRLr801BsRLwOw32f4Xt+EOWJwvL2GZ3KMFpmi5xMlZ2
9PXPBTyn6hf0LB05bJitNfg6ee90e4Mwr+9ICFPJuwI/kDsfWUMCf4r5tkTi9DB+nY0KW/icevaK
vOYz3XsL/lkIggUg3sa2NUMBEtbl4Z2mPFPK5eVC1wst2/aL979Dk/aENsQWWx37RHzptBSRRxbG
1UEX8Gk4mrtr8v+GZ92p2y5aY9AqqZ+FqNGtma3W24YWb4NKbdkRZDCQkcQFfp/Y0w/0mh+ZI6IA
36WyEXJ51KErKKUGrlp/tWcRsrCe/KayUSjZSgyWqJAaVajIEQsURHDmSck+rSKjHBKO0kPCRiLu
2chPqBN8c6dpAVV7/Ci2/xJlU+/E24jTg8cr4LduRXRq0AIR/SyE34vo8hVNqFOa8gskT1fnT4Yq
/VIdeLg3yonX6d1rKi3GcgFXXy0OAOiVUtPFd6TwojHpuCxqQwlHrtFtuS5WBdevODB39ozaOVZV
LmJTR5MKQx/I5UtfPbRHcoIVjg3jRHAnS4lz68lTNQx5VLcvmpqbhKgGECDUE+ohXkaOJAaZ0Kxw
lvsJV2PALNN2HDHEYI+uCrArMDp7VDL1v2bLPIywDXXPomgyt05osxAWpJ45Wx+7TniILMStSLJF
Bmt5+Ew8HdDyaAyXwzQujNMPe9cDA3HwPgyad1JMx0unvtUbb5dqWxbYmx1s7PvIzv1A7E0QDjFu
6vkASgU2O7n/DI3nFNsAtnvrRMmBFrgNfQHdj4UXAHmH7hDt74rewhIdUPoKtDJYilVJAAOtphSn
WjikCx2+L2AD9nyAFj9Z9Lmn1P/rPI7s/tElGiYlsrZFTYfRodaQKOF6n3bblk8b0LJTMPWJpMGU
6kkvYEj7cFicO+Ai960qU9GMZYc5VB9JLWJB+lpRXiD0ZOjqmG5Eb+dugIKq2Gz1mll+B3sWBkhb
wal5mtG9Rs8diHySzK6Abno5gltJHix29992tV4Z2mUWjiIZJxq9xCxGI06hB6uYm1cqFkjcg4UH
lokHuQ+2hmKOt/Drr3mdZf3QD8RoeL+hOdEo0fjILosYpsZpRzFM5JSed8tSYf0b2gz7LD0ongD1
Pi15QYlf0QJrvNE8nRkZPchHeiw4cyFeENF0RTUBl+KBwoby9cO/jVQGKftjr10AdjiQ93wqFAqJ
VBScN9h9U6W1Hy8sgS2/o9j1G07NFMILvV8Bvx4zvcFjGa3ZI2xhmKAqxrtbzDHwsdoOLFjV4nJB
0eJGkXMRpNbQiLgXhbFm+fZD5s82wk9/ChI50mxEW+xhecieOgHAjcltpEdJQlKZBzTl5Xjhh/pI
PbgHRVADE56k9XISX54d5kbYSb9okC7s1ag7RIjvfZFFYe2JKO8tbv6BQz2nCU2KVARrH744SI8S
M4kdEAnHCCNkGANENDKO5pRzaEw/bIf8cFslYoW5TCegDerRU7Rc7DPR8uzNXWG76HA3IraOBQt1
6tqauMK+2TxJxuPAA9pHIPFfciKDax9IP2c5kR1sex+IQmkDlmDDi5P9CydpQLuhSdgu2dWE8Swx
EHEZJ++I4KZSRplgmi5K/p4v3yXGkLHRqJiKLZrhytGylviFSPKqUZcj2DteLYE9Fskm27jH1lB3
3erxvjvCe4B59S6WrW+7ArnuLlHnLH4iii414AfMCJpGX9nDBPSxldaLDtiR0RM57daN+53QEJkY
e3GvdEpWorZ512+aF5DLoa4G1pxDox0tkVa/m3KrAl8F8/GfGy7e04ImNK4QvkLI6ytGnc2pVYhz
q73VOJiaxI8vbIf41SOntuiYLoB0/bpTxG/o5EYuBV+8l8hvqjM/NjhI1R8cUq5qwGsUV0uNJ3Cl
Lq2k9GhscRF2TxkIKtgziO4RAVussqgMx7dLtYEcl7L14cyqCdSlVT7T+IPPXgT19UdhyYlthQmQ
cRrUBxMPqRyprq4DJBh6dMH6BWs4mfQGxJ4LUZhX3HjF9BvbrXAQHLUB48x+GBP3Xian+8ADtLK0
DjyJHxCgw326SeHhre9bvc8Ov4VuYPhRJb8Un0m4lSnOoz6FxCWFe/8G+KZvEOrA/4z5wjGQ0TT7
kU7dRvtw0Rmag1KI+vqmXMAUG9OfBlmRbwhvX0WbgSwOZHaFdNK28VCoRyyjEEJRKrjQOn5Y0DFa
r3O9Aw0IRthsmhPS8qXduN1XDnanFe7WD/Xxwr0o+kc2QGtLAEcsJh5N+kvr+wVaNVfggrd1rfIg
PlJTAAO9+L4xmy7zvXtB1nvOImAspY5oaEpW1koesuiZnRh+BglMcNAkpTB2xmSQ7Yb0zxDJXr8E
2xW4bQqYSMUMMjtIM+OPzVUGX9AecMxgF1ppqM2D3JG2GaGc1TvrwwY4+dg+sE0bdRsAHBo9ay0M
X8fzLQnSU3mMuzS0/MqBdviYoaHvNn97VW7AjENCHFNjFDw68eBxx8Rn5S5BLke/KSpWMtNLFngq
m3Wt1+bHhJQQ6KTvvzZOzzTeo34OD/dVGA6PhtPsYyw3NSW4Jm/A0WYjEOp7m6a3cehVWum601Ha
1L05jlKK4/iVsx5/fwTV1FXHzDckbs+pn6ugjMBe0ZH7nupXPM4fOcywWsC19809Bz8lNLtAh8tV
AW6TQFf7VEWLxkM9iq120vG86pY6o9ixksnDD4JdkeorXwIJtYy5lhUrYi4lR0TfJoQOKOlB0D4G
UT5RM5sDT8UHtWkGKd3YewGMjYI56jxtZvkLQETBrrdXACK8blelZxX74+wRzNqxRxqREq7jQLup
xh/6h5ms8g+2v4Xn25ybIHF4twDL6ePxi3Gp6yWOuj8syGrOu8G+CDUkTxwpxbxxWnpeTb+qfZjE
+hlg0rFNsNMci4ToZDKRrq+aUPU9yeg/gSVZZCixi+Pg0MqQKhIhZePpkuAgc/IYoyjAh136ty/P
pgt1mvG2TIbe2VHt1/SEZPJ2+ZezNPNvvPcV8YVIbZsL2ge8K0s1Bv6cvgGheCDrXGPuCxIxtsZX
S7qN8xCfYje/uZzDsN03zXB5dsNeq4KbBBDNopujdLOhImVmiPcjn0HTK8D7rrCpEOrXE7LznSNh
+oIrVlBVRzQwNW7hlrwzkbd/kV8cd35JvNttXB35TsmsyTn+a+VxRhBxo6EP9k5AFTk0aVCrjvHF
jrGakiCBBBFWBM/v0hzlgBo7z13MDB4NjC86xIIaH+xBQCjPyLzj7Px/UHu6t1T3Mf6/xJvpnXvT
0MNFybpuMbHztV3rzA4oidAT1VY9OehwP7hC7ASAmOO0kud8mnJTlgYW4IDZF0vcZpbdMFdENFc4
mh3qE/zgK3ToBL83sj+4w8a9EJDB+zF7Ek6id7aTa3QZb/IwU1cpjEe4dCBRjs2EMPNyM7HBIMVp
I1mOmy5nz0/g2bxbNBd6ERbXagE2p8oNBnL8plGA16PLDd9u4cWhGt5wOk7kjpFGIKlzC/OCrcvV
dxz2kWyuJ6qr/LfRFK4wtwjfzo1FSKIQxXYfQ+jgOGEsJ+LB3Mw+n/d1YmUfWbXRROGBHyYrXsng
8pA6/P2b9GzeJ1D94KcoU5T815f9JJ086p5Zw8j8S9xUDVEucr2LAkXwOkfAgyFSIVE0TJm3joPu
WdyzY9jj3HPb9jv55PmRBxb1lgxEuzXGPonObPqTAUgsKuqt2+0JCkoHvzCc5XtB9EpDBOi3U94n
eyXELkjU7F7dIGtKMnRY6mhVy+aNyUrP9dlDfC/sE5rByk22tG3QL5m5zsQdsniHb/F/rWT/QYtS
grod+e1xdr01c2ILHLKDJeY/zk/lnFFwRFJXZUxeU888UCVy6l4O/yhYPfIwvr8JYPQrWyUxSQgU
PoUHogTFhlqss6y2oXwLheGStcXPO6XGqNSf29YxaArajOiU2wrv7aJDXM+YeTSGg4sgp1QHTEGT
ozXd26fY/aho4z/khC0VhaK3nanxS6j5XuDxs8Zl94413GblKJks63z8/RYpa4UMdIPol7IaeexS
r3RlW4AEKLQXQ5FTQ+3FtLBbYYscFZOpWMNERV7/ozpUJQ8cYo0ox8YgX9bl3ht5FcLqJyr+JRZY
TwqTJ4ZkZhM8WBX6F9duBwtgU28kox0pFt/7b9+VbHs61G9uR4W2XmAAiaqHfaFmfhcuuSEEyOvK
Tc4IaMQqE7HggW8OBFpbn7cy+aH1SP1iXi69lYmvIvH/TxJHNYwKuOpoMyyoewNAtpI1qMz3tyqi
D071fhWYasFCjfazxfaLYGLl9mZo6aLipFcPtgHN+DUzCa6wh5/ppK7orISCp1xlbOR5wPLsbvss
uGf6Uoe8ks70yeiizxQy392nyKFlOnXTnzEka4ZFdoGWPhT3qTOGZN188MK7c6YXqLdm3X32JNex
oXx9tLPe05gWG/0nMufYDqYxEJtkEMA6Dw/U+l2boBvF9+4rEG1Ed6ZTa6zLbGNnSpkt3mB/BD6N
Zm2OUysoHmONrARYVToiQLYTaguiiFhU5SD0TA0Wct6wmrANnYHnUj7oua4PQ/3M8U2osSQlxIsl
iG+4pgnf4yKpRgSwzNEVwtl1rypZ+VfmIVdcvYFeWDBHuonYWVUP+GCGUfMkIUArjcGlV0hCzGee
xUhM9qg2s2SQUjT/Cr/qn6/2vjmZfHcgOVByjlZZjr4aiQdM/aL5eZSIrtUnfxA/ip3VZQ5BWbdl
vdIgMdp5epC8nFvZRdTvucvpEeAS75R0SY/pXhvlrS7rACrKV0O7aWFD/rE0BcqPhoXZkzYgVRsU
ZKQ2xzF1Z+ViHAKfBAQC/UWYf5ghhHRn/k8l5xAbPDd7D1CHMnZUcPzjUzpKJWf3UIiw0ddDpFt+
XWmTLoNIzl52HrGf94dBBah4+pX7KVdlvnwpRRoNAgV3LucZlUvX14OgGcamFnUmn2Wxp/zkjpCg
sfhxtEshIF8NyEtO8aPjRaoJ3yIg69hbFW6uFwo3aJA3dUlYaEcZ+LVEiPVMY6Zeky58mzLqKBNi
kmwf0qAgIN8Wni4UtH2coGSJVZTYytnjbc6TqdDoRyHO5gaFezRSE1U6CbY41NsXLP0ZjTRtMBDt
2E42ZCP4Qg7VSFBu1NaNJnIgzARaW97MwHb0pUUJmMkOGayY/pp0WcctmDVErbIx9z2SgX6RCuMR
b+y5aaNyKN/OPT9sEevU5LBMbwn2iqx6ZUsmpiOAOso7lX+H7BE6FLWlEKYqBrMnke3HGzTUDBpS
8+9Y1f2rcstxFi6L6w85qCIG/CNf4oPNddlJ9BK/WbO0XW+QzUfGmlWr4YRCHFfMJKf88w60V5tW
sPfb7gsX6VvHGmKebisz3B3xuq7ocgkMXQp7nK35BGwFx4rfe4+GrZVPDJKhfPbBzVeizUkJzLgX
bM4etwA9bVt97ZzdTEPEOg1hV02gxfGSrLZVmHRvFQmC7y7+Cqll981hT6voif/N8Bi+/7oAeX9O
wC6nCSKRuFdpMYU6Ia9iaGpLDTqeku/bIsdLCaiy/Wd5dUMHPjND2FrPt5yuD5gzC8ADZXFX42wa
JwyusVkEID+EEvbvYeXUeP1vOymRGh76RFchsfkEkQlcCfedudGZ9iZCKA54O3/GDsdaF/LNVNfK
vsnlm0ZK3AWoeXWslpGOpBSh/OR2kEJhJCF/79XEwn9tTviqIchhKz/4lOD0qVnZclIv3+JfvXWV
iWAegTPtm0fdWaRvIIiT1WvJo/s3AwoiVaiz4TE7TfItI/iMqrB4crIWBtPgrRv+N+mDW6jMdpFL
FPakam6JPYelEoWyUaMi2ijkCo0lzTJsVWA+okornJGBvpWD1JjPtFnEt9OEncj85a/e+eXlKlkA
/rl79ZnQ72toLV+lxE2n81ewGKT5sDOGPOa0/8xGtn+6E873vkh42xVmkgCbN9sHcR4FBo4iL07F
cAw3qal5rssM2OWx0Ym1gV++hIUq8NDzVr3APLkGejYVqplFfftOpSFIba+BMKQSf6HlgZV8HKwY
gIl+/nITIWeH33Iz8B+PiSX9nv0+Egj4ctmb0TVycv7lKwzGm7KnlM4FX5o1xOjkG6WhCTjJcCNj
GZXFnFb/LeLktVkFIsNXwdPl7fr5R7LXRbFqlF838oCqbsw9vTuNBgWUDU6I1FgHEEEgnRRjhPnY
LPXHcDBHlqRJ89hiRJrOXxfNFWBiMdHk55/VUaumxee0VpelpjQk85wsl22y+H6L3MkL/vV/T07n
KBAWXoJbEAFnZ/YiMpTJfc90M/ZtYie+p7F1lVUYBAm/Z98JfliEodvSJ/kjCMgVqS9k7sLUEzmL
+HIjYOZWCAfVEhjsRDAFCBeePJCSmBqam+bBabcfiz1t/9ro/yGym/BSQRgVdHC7Ky29h4O3pCeY
32RfXuTvHQVIfgsbCc+OYz2EdvQf+kcpnzylepWDvMzNqRBShOcAUqyYC1hSMZ7cI8GEuKuBTM3b
dwiMnZInsp1HglvKuQtagcK+zlmF777ofeo2SFs1eHG9XLo+IhC7AqrkQP3mvYh8Oabjc0G3AVLo
pojY8Po2lPBxqZbIsaFske1rAykunE46YggCr6cMJfX5H5R3y7YlhDOJEb07IblxJrJT7ERLR9R/
cxcjXiiVv0hAleEZZCBmP+Tu/ckRlAb+mW3zyrcKZPGKXJchJFhzlXJnjzFM7vBDy5tEcfX3dLbJ
QwmeYld7+0FaHJ52BgRXSFrwr9rSV/Z0moJrj2tBG69O4ydbniKvEnFVk/nuPJtHAlbD3UPi6OTk
zv3ciHtKLfHn89L4/tnqzAVB8DDqu4Qmz4hReEq621y6fxHiCaG7i3SeAouYAWakMFCIZFaY5Wgh
ZFFnGlO3AzuPPDOCbbuoLc92Y4gJAwlx5ch0iz7Y3q/e+KwV6U9jX22yDkvLRNS/1zQi8yHF8lcQ
Ikj7sL3aG2mtiZ+QwKiLQs60Y3JC3YgLfi5enIral1RpEf3DEC4Wgn8JpBq/1XHq4Yu/HYND2Lp3
CE8LYsJlamdWpsuxa7O0C9aD24fHaPIEg60Y93AYo0nHOdKSCQ3hFP7dZOn1aN1rG3+JOHynuWnp
hOyqro3Ucf2wMryWZritItZKvplQ8EJTL55DXchzLE3WB+iCyqtk+mnRqjBzFAdOwPfD0TFcjuoS
87D9//T1vC5Nl8jnRyle1rxTVqUHbwRsvv7M67txCjhoNqMwRYGBYrMuLFdacu2YRbWpaVVbIXQf
SA1b4zgUFZ2Ybz3MaDjKsOC8asRZ+/8UZStv1bUbEVSBWP8AkLpm14ja4dlFqlmLYfMED2ekOlYd
CtYyF6azhVhImIeIuZ0rdfagdOp63vGKg4qCBpLTesXsoV4878w9CWLh4ezECMB6wfrnm205fFz6
aJ0lOcAfToP3LrePX09XJ+RcwiRuET/upsn7LFJeK04IIqqnuZpil4IRcdT7vMLDn7JTCQRJa6KC
3DnR5OazhsatOEDXR0ICd4ke8gjQ1jtQZo/MA84Bh18dDU5xsaamV4dUr4kk9799mKK5qKPC/hHn
5TYIXWVu+nwEvELaWF8DJjZSreiBw4eqTbFC+Vo3JyQNuirMOSTKzg3eFIhoOqdg9pLJ85Jd33VS
iUN7nlZCefg9bN2eTRLIYGAeO+N3JbH9Ix9Q/FDDLAIWoTIJ9UBVzx7ukScueyb6/K7x7Vz1bBEf
7S1rwCOZ0UXhcqLJ1oYavvGCENCRd+uyAENOwXLWadSeUrP4Y/q/qfR4RiwxbBvs/UNuPAtKdzjz
AluZGeYThkkCfL6JDMqlBX/H5sddLaCAvjc9idQl2BKbrTRQ4R7uQs2XybvcxztcE/bJYYX82f5K
JV5PeghPXzVavxax4gUxFblc3QBbBopyD+6elJI+aLpymOX0OpYCmjdtEUxxKxdfYoDJeWpYjb99
TCNq3lwngLmr1j5zV2zZlQOnf99MenHfCcH/4gLvJWwVDYXIgqYjPToJJsFk3vs57pZ3IL4eByx1
WVOhpQ51OvZExD61uIGk3g1lqAoFXYivX8KUogwf7fKTL9TUD5wcoxQH45mW5BO3PNtJkXFisG7m
Y9EypveLpNjxGzI9g3xOu7u2sprc4pXCE//53/g9UK8T1X7Weqs3B2MQzKgm5J58pMgjufxsQxfj
P2SNbyUOehZDltxekKMaPALFIVpK00zzo7tRg9AWgBuJ0NPECT/ucKZKlsOwHtmQ8OpR/8hGwSCI
gAzQFd1u4/JhM6m25zHPU52rXA/ydsctwBQEu2qbQKlluFVdthXWrG9XAq1fQGN6qQ+vh0FuDH/0
0bgninN9CDQVeyI9wkYVPS8pun/CVJqiEdTABwmEphb9bB0VaShIpHtqv3t4Nu4z7HsxtA8uSaoL
Iz/KkGBkUOgZblQsX3TOxTNRIuXJBnggR0OrQv9N9mXfNkawyeKAfE6LAuGzNmlCbNUDcC2zYZkc
l5MoYaU4sULgAPrHGuPVKV+bNS7Ndh0OYKOTRQe//OlX/NdaVGqbk6QE0ODW3UqQC8XBUu4vYssf
5bOIUoVNVD/5ZMcxMiFVYpz1ADsoqfDh1AffhhwZRzLYo8lOm+BbCU5d3CmY41aR48sa268XiwPT
SlgGNTZePBxJid91aWjb5sVS5Bc6deemOuy3u5WKZhnpdZCMYUc0wO7KdQIVzfo7n6nXWDPUV0wT
oQgvo/kpL62PFQZ+qo26488IkpS3fBq4qa9q4jSUpoLzuNiRwNrV0RSx0CxenlPr53XLHGT+W9lS
MBaUCrver24RJ4oemFA8gQPySZeoiJ4u2kwGTa1W9IyrKK3LoR2ux1jZXf5JpFIhCIkOlngQ/EyT
ij6cj7QzgDASME+NA1lczHE/LcGlo8GEyS9g/C9xVDTajhgNLFYicwfPyQQaWPvPvMXCQmXXVEko
Iwq4Yl2cEPqtp2/S62YrFlpyKq3F6r5qW3HM2pMn/OM8505LlnSSnpcanvbWgWcaj9w0WGZX0LRm
h2jS8bv4KIOLo9fb3kBOYbl+XN5mVaTjHApppFHO8rVDviK8wDoZwebu+H0obakL8Zyze1hK+CnZ
R1YzdsrA3wz32Qeisg99JEslJvIiCM58pA0E2Hlpx0vvxJzJ7qE+jQoOsrEceBqnnc8DIBnVrV//
0yiSjNcc6TYg53TYWprhdLB3v73Kyh/1MXvuWan72plh+Sd5CRGD1thYl4qaO2SoXf8vv7dYRUXo
28JpEr1T7gVc+vnCY7htV3d1Qmag5xlUZmz8QbbaF3oUKDL0oB8+Op6qr9fBKrMYPHusuoaZuc6G
xqEbdlnJjJ8odDr5M45Pi6PLcEc6uc6VYQ2lOQWUCI34N4GkmdkdgLeEw/fQXZI75AKLTFtZjXB/
mAe4OOFUrltjgDkWOVa2a1uqf1VBIku+/o+c+a0dKcbBXJ6Z7OtdBqle5iq9tNvhKWyCSai5C/cF
UzNef7nrtAgNE+a4vFzrPxxmyp6/9JsEPxJuAEXIJm+GiyXflVbOuxRdsJlGgK2/VqUm1/omwDnd
kcQ1zrAqiYG7uohVvUenKdd5XclXYhLJ873kxuDz3g1BQXITGKqrFGZWVBJZ8uRYj2n78wYjsaXd
7bp/I9L3fjT5zxCdJ1W5oCgaQglJkxgOJ7Zqzyzkxszg6jEeP8kbfQz/kyuxwLIrFdkNsxqGJoBE
fDgMAEZVdc/MfpXXdMUooblBMThHqMp1GnonolYVGfX7CMDTc35jRfgUOHASLAOVvWCgG+t1IBjD
Mi6CCnwkyQyNHmSmSLK1rjC5D5cpTZwIF8bRx8Vz3ycWzyTq/XUjGRzxzi+Sij7GCrz4bYAabvIT
BmX3fAnrNI6uenzu5hg5SN0DEBNjjexouIkO8s7IXFkASb2RKyNbfEYkCdzNnBCYj8DVua0QDj/g
e5awC4uVJS1iRqF2mlYN4qHoPPNcJs1FZao9raM100DeKghAsoXBh8qKOX23fSw4HrT5gNitsDqS
bJY7Bun6+/HeKzA7Pk3/91ndt2YkFb+k7d5Fyedb1RuDjm2+7vNtAvFavbtlHr5HyowoUJK40PDW
SKrlNjTZZgxXd5ObMrQRgi8KD2RgrXAzKFc4vspqdeExpXKJ5MWK6VNj+Qf+skb09DkNM0Zy6nmR
tIuvj5c1nKruCWwKQAZ8K2kSEamIymFFoa28ypBGsI9oJIq4EgzDTjr9FQoAjjZ/eZg3lxNRdmYV
vBfv4LGD41tAp8ykJalYJOePCadzSR51LdHM7daNHrd6lEWIP4ePKoRsMptudFz05lwPUlY6Funs
j81evGWQodd8cQ9u9PEQenGpX1m2JbD5lKupMJwQj+62z85Hhm1ju/ce4/0RlInUSRRLvTWJPjgr
MDru4m5XeV0hCkvY2wi0QWE1kWetxaJk7txREnxmly7/PaQuDzJzfge6vNig7M3DwaxoM+nFToTs
tIa7HVtf9qBetjGVAY2Yh/b5f0wMaT84Bc1ZRjirAa0LRAizZVhkvTNxy/00mCSPcztleinNiiwE
jqK9h46Z0+wHGsyL1g8RGLu/Kihdjd7z+XxfkVJ8ylUfcbwDMQpY5PWy/tpttagl2MstcdOSa3SL
rI5TO/KUyyNe85oZWTqYaj8byIRGxQquSpKus7EiUu9Uz0MMxZFWZdAg9zcGwGSpEaPe3B9fWqbj
Iv3FxVTg//Q8x3+rSf7lVyAN3pZghbmzP2Z2ie2AGxtJVz0IwPGGQAc6pCE6KxzzrTJ3JpgOtKM3
NEE0IiRyWPF+3vhl1GCFu+TQem8aLt+ocJeu9uFjfBK9ji87AmMNOWYOzrpoM+vp2PNf+Df4tRdr
uyJPXQjXtM1PctlIK7NKLPuXG8QyOePSc8kRIyjkswCYNAByXO3TMuUJIUrLVpQ+AFHykEbw6I5E
4zp5KDdHClXf3ZPRqklbCa1cvqu64G1djbigeLzY+hZV8UYo/EAPVax86V9x2GD1tIxIC9Hm2wO+
3fDfWh/nSMa5jqdMXqBe5SGHctDBRfljEXmYeBFuamVEOpHqHdr88PpHse+Dg/4zwj1kfPEWkmEk
H4F/Lneppdf233H5Jx7b/FZ4Q0OLOi4bLTyj1vAfGPnIOum4ELEb0ZcEChS/aIMYDl3qz1uf56IV
Ebj6lPson/Y/vd9Vk7lE8elgtcvtSmXVOHkFlYlwuv2NHOnyEyvmSjTLs0GkW657Na0BOuwCJN5M
0BsmtDM3ft85wylMOHdvFzrngxFKEQqBfbRIyPIFWN7J94W6tj5yFM/VgEuCtg9CmgNaQwmfK8SP
7WvgGuW77DPlC/IFOg7aQWeGg5vAHfATjzGgrFQRGYePwS2FL2JI0YIDu6EWVqR1G4ZfWPBpWoJO
YS8rLMDqpt7fYS/hjW8O4X2fhGEFI0m7+TMM/GyBp8Ty60t5GHI0zjE94LPw1W9KNyX15t01iIo6
06/pu/JeYIGIJpj319kGMXjFFiWo7tPvlQNL+j+xGjKt6RQZJUB/u5mWU3qlH8PyAkNxG8cihvNa
WBr12/+5i1UtUE8/Y3NvDBb+IbCNKgKyxFymRGd9epamtnJeC9h0eMN2tqSrELC8zv4NSAKRIn2t
FZUM/3TCe4rBocgoGQdWChETLkpICr2/9POC6DJ1zmhKGGdiHmgHZlf/g+4FfS+OuSIb9tPQFlMT
KJubWpFyoO9W8psmwMIlz0imDqTdTNU2MuAWJe2f6HCcYMQH+523Vw+BHJs7tLwKN+BDtEaYcdsf
44YzjWDreI9THz1WlQtj/aryz/hEWeUH9S3DfwokWnECR0NK3I9arMAqa9+3yv9ZcHCwMZ3iyLdO
OgmuLjGqeee9Qa7c1Y9FelLia2UZqPGgv/sR5kyvvFeGdV4cQbikBvpgCVo5FrNEpCbY7iz+1dwg
Zt4LoVJsAb37xN2KEC5PkGI0DTGz+NZwXYAqPkoz5So08KziQd7aa54Yq2Z1XU+DtGmSXb/BICwD
RW5KfbCYimclqN5gbviRAQT6luw7arpA2yQBMyfMXCLNRanxE73e78scWvlbXmsc13og9WuZP66U
91PEUAY1bUvQDZ9zBfDIt8RkLwC+lED/T+4drN/4hH2mcphsjnhUIioyS/maImG4QjDXvfk0mppt
qdVcJdYtd8vM8YiRpBKJB3ycMXNXrtkBwAcsth0VMNtMK2AUrcrroj3My1BH0t0b6Hn8Syf4gF1J
tnRWFAOHxQ16C6Io0LJjyM9RnlAYw2clCQVBGuOhmhU+GL9DGoNhh8v6VEXDMunFGWIODIBO0Igq
hTB5p4UoGvi6FBmTWbhM3AqRua4p6xQ9smyyQyNBPiLeibi8KOfQTKLCyI9tJNeyOC+v4S834CB1
cUotbfxhy7i3nXfYVFEhhAlMOTlT3czzZiRnTR9gJeX+bo8sf3O3M4Cp8ttb28E52hb7O3JYNboe
ehWWu3FJ9JLp71QYjm5MsP7g0NUbfoftV3GeNo+PnPAnEGary55InWkCXArp6GofK86muAeeMRTG
rmA9pCzw3s7ojrH1/w+vFmazQESWBSWDhskE41pwSRoRw8KnKF3uLcY5utdQD+iTthaiR5YnGFYW
ETycaOetNVNupDM+BKqcIAm88CcOjEpldIse4FknIq2yl1rHALNjBD/PBGWZZgN5fJ9tHMzsxWRM
63zurLcBQ+XRWWJA52vpW7R926fGR41ACilxSKQsZkW+6D1bf0/g3ezXu3XwOFGF+7PdHIthLWsz
298r+ZggnDPzx5lzC11wGw5MpJ/CmZgrYLRYBLXSB/TxjowIRxttmQFB5UZvhERsmTFJ7ABlIqI+
WgdNFDwm7CmlZBnktp9YYxd9OBBU84F8yX+178QRLTFDJTNaSQ8tjOc425HgyjWuJsAKW5sK6yht
7thuekW97rseLoqv8AeIW5maoNZ/BCjajz/uhPQh0d/hQt3LcoxiS5ftq+0v3iZRT1c/gNO+6Wpm
wRddwfQNQzzK6x9w/v2aRr6MJo0IyIwoWsld2AICfBrwZVdQ6a2zlO9UNHE3UXfEZEEiqLXcp4jb
kYqFOaDNOylmelZkk495w6nqxz9yV7MwOZmjQWI+yWr7xJw7gjl+06zpuvcO2N1NEyos+EZxFUKo
ih1cMQbwIDV1GVId4cyAjkpMxdCaQxIraGpguhZGNmkVjW3cifOAZYFgWVy3XgW6NluFgnnoLJiD
YLHNU9l/Y5IfOfoikmpszFzHmuWAzfdHRTudjAcn0awqoheE47g0VoJbFxe5krfuf0cx5nyN0dpl
acpxmvOh14TXqRqB2WZz7Iophr8xgLPcOVrAC5cS+fw0HxdrCVmu/DaJVAs3TntVhrp/qe6j7aqO
lqAvFw1DbHbBGWvXQFwjMkdlIG6es3CFAA+2ZOlftZP7sBxpNNFTiUq0LQm98bHWxcZgrlb1fdn3
sQwMxsEVFUDWiwVJx42H4QC9wD1hqpXu4aUlZ3ItprBWjKgAWto7oHAvoY8Nct17HSFAMKX27G3C
j1NmolHFNpRdDlKjlbGjzOwr5aITbNNTx3PBCumowF4FPE0/KhAlJzM+iRbxXqE3znuKZzCj+1vO
53MBTaFCYmfnq5yBPIOMltAW3FtVTdBaI2P1v67A9CHcH4+SD+E/fNbayvYx7RPisCki30l5cfiS
iCfRt5USSf+u9Tj5dLsOSSsfvRKIbjTc35Eb6Kj6X6GChVnUgS3LVsLvWMUjIUOhFBXp6To1SGGF
jXQ+fF4TO3FKf729Wi4b/E4FTn8WJ2pujFny6bRkU9gWiWceuEM8RFms6z1Tn4nKzWTIfmz3Fav5
UlXlc5gu2h1Ls9IgfepztcEtOBFKod4FN3Phs9oCcnQ9a9pHT38XO00wEiv0Yslv7JivLSq5gb/W
6x572+7YxRpP/f2zfGfZyLSM4tMj5iprNMOUlLwZNtqNAZdYzMHSfugwadSw4idsnoGuSo7WI9n4
lAw6rMVaMUOnag/aTUapD5kvUCf2V06aPfAkieCiE7muz4glGnfpS236vFFqfmQDRtnh/5NoIyjs
06a1v9yHOkDmDSg92bKekhXskBWNzFMHZV2AIJL0OtP5W1EaMLp2aXQGtyphn3cbf715jbnlDfS0
iehapxkBsXV8OALSthm9gLL/aBCKLZf0aREeMFLTTDZyF4FMCDEqD/UGq/LB3peYN78305q+OpiE
CuaEYQR97X6mLZr6kvYzUV2q6Qy+niH7KxUFYJ8utQ89M4agmerdKIs0ZlcaTEvfhvaGxqEhTYW3
lfUvKVY7tUo6FM3hAaEZiJYWzF3+99vWQAYAJP8J6WHp4i2WBG+RUgO2awyxbYjqWnbJ/03Cg/Wc
ZI9+GJhv9g34yUmovuphwr9bi/qdaocb9djW4zkb3FDchX9RSH1LCt7ybfsJyIPyriDIRiAqPdlZ
as0eOss9TtT/+150BYy6O2hm4AMjiwJ4DJGLzDjdxnj92A78FxbhXjcas03XCGAIhHpHBmyDzLAc
MYaE3xiQ8YbEJ8wDeOEoBWZ+BoC5kr7qz3iKzzRxZN9P9MZAq4/qc9Fnjz6/MCml1tOcVCi8lcAn
oej9R4z+6UtEulSjujjE+6xi0VLJzTxh08u2aTn7op9u/9Hz7yycXSmJh1/1p5OL9/Jtdp//kS9K
fciDfYnnJTBNCVclY8f3zFN2kENSAlOW0FwlfFX7KfUg9/RAvI0N1LWRz9myPIazMFZN7oMUDZki
N6qBpR22WOiN6o0eIsRaTUp6y2jHwgK2KAUMjeNzB0yUQOnrDYXnJgGl4bCgCrMUDqVnJE2ornaa
cP5if7szUJchcciOVhlWYGiCNgdhHG9av1w5DJNgETDIs0E9ApmT/doENpLWhPjeb5j2NDrgT2bR
5vhy6CF5XmXjhCTxe4drJVDUhqophft+w02CnjLQizfvLMHZwQnN99P3Oo7bD86qkGEX4qzxKhaX
B0zDv4IdHDXfqAIaVmU62/YanfAQNAtgBEjZu5vqaizmcTO5H2KdtCYycFEExevP/3MCW/JMq9wh
5egOLchR/BhUFcgLhMqvqJFsVq0BvP/2eXfP6pi5N8BzWOMmaMQFycukK/cGA8ljIlSDA2eyP9JQ
F/wOFwr3mJ70IlCu00C/k+/amsVwXIY79ukvXJ0DAXxPZtcbGmQCT3BDKf6G05ogR4tDLBYdR6Rj
/RJThrbkhMVci8fkacgYfU8x9sfkGkLbwuOjqhCRAqiRQmMLdirW5k2noJ4jTSk9CPv+jhHjRwWT
nVYJKtxlXmhF7E21C7q/SzNJJw+xy9ePOI+2u2Karp8Fwu8jmKc7wyMK+DAHEFwlxcA613SuUBPN
uKUeYTssgUJpTyrC9Pm3wnxi1TAsyvpFlJIBberzT4VOjYldzQpSogDNUN0AR1F+HiwA7jxtJNIU
T0cTwe6TqHzMG3yehsBN6C2Sml6XXlbn
`protect end_protected
