`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pVSB1fdp0d8mtg3LHrLYCqADYNQv1kYsGBMv/+K08aLxh/NLENzMM7hXXYld+2Mgd7vecGpdaC3k
gwoJ87eJgg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TrvLQEi/uJPAZXHsPaV57yoJ9EtvRVNbWErIxN3rJpRzIiClrcH6SWry1U/juttM6Ef9Hp5zSiEl
xNpXxoS8wD1iGQC3wTWm6onL4lbs5dCr5r6SHKI+yRvk7PM0lNGSuxzJxiESo15OD+VI4TBDw4Zt
hcxOQOC9HXnv4RekyhM=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g55PFOQz5gBNNuoAKJA6LG+Go3evy8K7bR71fr18lbAHBy6BXY5cxyMVmR6iMXA9xjvLNX9ZwFxL
yW9jhdIKz+0phA20qrgB9zIyJLsPj7lBLFXWAKf8rmqv2GMRf7GqCtYK5Pqn6bxMwn+n8j50ca2O
X49Iq1oj34Zh+mics+4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JjYKvrh9MOLSA4mR//LjTlBGaa8xCFhn+/gMizL6ZibhVKAfMan42h7Ih/5YTGi++UTn0LHd9NL2
NaEQm2v4o2/CYXMF02K83EGT2I0yUSTUGc3tcxpNAxg390x/Pf1S4xXOwpqZAYLjhWse/4qzYHFe
iIQp1rnWICwKmFo+ZDG7yZ46pqq5zbSoc4y2p8g2Be/9TN+Y61xI7+D+EAu7QTdwsL8a3QMsB7Zo
r8bdBBswbfd/oqL9KLKL/Se74397O2HGv16SR7618OwhGC/PJGF62sCa/WzAZbXDjbk7bTLUCyoY
71dLV9qD6596pGntd7mPSMKPXsrBqm2dF4MJ1A==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SSijEQc3z4IgPRpOXyZNPGTBKNNDh8UIUp6Jc6nCd2BhqaRyKvYRVaSbO28FxPLannTOttVNc7kk
nl077g777DPyzXTsDcYVVSgCq66KzFzd9air6Rm4YQEnULnroQEEBvsGlrlRApzIY13fCR8Q8Fes
8flh0wIvt1IUA60/FMM3YwNPai5m3k19RaY/qsBdtTNLM+8XqaS0XCHWnyA2QHtb6iqRTQyHXNpO
tBGXOMyVMkyGUq2FAx9nYlTvIbXYYvrUtsQaGxetWks9vlDulbTRAnCFb7GU0+h3l3y+hF4Wzkn2
o2p95CyRx1FQ/Rn0oxBn++Rtk6p7bYPQS42cSQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L337KT5q53NKw85qdeX1tBHCmb9rh0WndWsKzAyylJ7jXE+LkDsZ1dyUX2YUpfCn9BKLEH2MzATq
tqzbaiVWOu/xeMRiU5/wkXL4qEX/dKjPRSJlNBWwDa9lFGbdFy89cWFoNvS+Teu59m5yiiDnIsEO
MXDu8nBP5UasM+BEuesC1UlPIu7vinDhIbxmSZZQfdQoxRJrJhS5MUcMYRs6Q8mNJvPXbo1WhUGq
lCkeJ1Mwf+GUzVwd087Tb7Hf3TsU6tjTfAyqJFoofzOBAnyD237xgkHu2B+/4AT6bby5CbEp5ISZ
1Crn+G5ARbRRqoqaFdx72snFnkZFJIffkdR3DQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6128)
`protect data_block
3U+9z3xqvHNIcHJ4qx56r6NXAFA3iXsWzTxZtyMTPdrGx5tKrEnHB10flD8IZCSrwT84nKtML1yh
OMCSeU711Eum2qCVkKVhGiZVj5RpeclNwJMBai3jK+5YpyRiOkim9ntZ3hmuu6XMbdCeCR7wYe1A
r9bE7kD9zSPlUH0FBzsoZY3qkRiVajja9BiMjJEEbTLM/wW1zZnvYuC+vpGmHfe5IuWthoprCYGk
SfOICXJIJVkGc4IwR/bJRutTEnB9MBh1HaI6CocikTOrgbQ2jVyk1Q5rQOqi7WZD6kBkwB2VQZZv
jqee8XcRnJ6nY3C9mA7udZQEuSxX5ZCWxELqd1O5yD/o5NMkpgv20sJBw3bx64wPhkuE30xBhSLu
sw+QFZzeDYUPCLQXvo3ehqPBAKJCbzehqm3KoVa3yKgL42OZTG286QPburTF3yx7VvXFOf4H/4MA
6Arh1eIO/k1v2+nr4T792yGfbmfUOSSLmqm2YfoD26PUY/7+GpmJSdeprKCzlVdmDZarSmh5Oi3e
ZWqamWKubymS3wVpdqzmE7leGVbL8uY/LU43qjMmjTDtv67wbBhb2wuvaLNQL55Vr66hsw/7uy/7
yNekerY7iayt5hNhbf67hwcDRjT6yAKbP5K6zZO+mWd8xay9mrDNTlIIhe39aFeMJMrNtLKfBnhA
TEPlm0cM91uBkbwmhxiEcet/fuJOEJCl3+HEZdDhc9Q/TICyShFFKNtY7d3qpt6k6xPFCIReW7O1
iPedYTVoeAe1UWFjBJH+ae5odib1E8BITFFawhfCzmJFSrhWAm82u/8WEsI7sfPRaC9UEBzKo+ku
BAUbOyYMK/JU+8ZZ2nSNOd3iytX4RqVkWROYMACmPW+2gnJax2saO4/zwuKjWgsx5OhZs0i7NQX4
4L8+wwqq3xzeFZdYrPHi1ROHdfrVPifCpEcIOc+uswCgVgbw3EkKg5nOW3V5BKOHWkN94msKSgeG
uyS1HxCYDeNdRuAPCl0j6bMpL84B0XTj4GQljbGlaqP2yCe/gIUx7sElI6TbNB5b8xxMqLpl63rl
EPB2SGlMkMB182LU/f1fP0Yw8gaHi+sckWmkQq4FxhhFyQd9nyvrvl9206dmXd36TOr2vRuHaB2O
oaI16x7HtnS9JXKt8VhMoGwhLrOZVB8rLSJUO2LjkF/QBroKNVuUwZaSsZWWuSus0JaXdeXsXbda
y5XE4RZ+WMCMm7pjCEsXulYQdF+8rmN2M/Qss5ayRRSM30fhjelOzBnHo8nPFsHV+wfrBgIG7UbO
xMzga2xaqG7jWNSH9RiMLOsvgs4bPvRCFQI89k2lkWrHxmr3VSHOk6t+/V8Km0T0qCe4g3HdEWm5
w2lvi3amMGpOG7FJRefTiwMHHzY3r3dCdc8JxWB07qpnkOETZpnckHym8Dqvsxw/HOhG/iDtVWUL
lk0X5gvAe12NZzTK/1KhHApUUMazqUElgq5rScqfS0085j881NLhO3aPtlfDryKgujpXjIPB/Gyc
Pe/7xuH5mBxBniEk2WZtnuIMreQdFl0wAkvL9WcVtCL9EmKxW4sc6HQ689HdMo8kQ4khgbC4uEls
RKEIxLHUAvYnLp0eu3nT6aqz0Z06PTTu1V/fv6F1gE/CXCH3ESvCWdngVZdE7LHx/d9lhnFb2Asv
lKCK/zGBB4JyjHY6eE+vnTLfE2JM/pai/YqgIjkKZB3VHUfbxYeItcLfIK3zl8j/cPF9o5wP9YrG
YFxCxPfuREyFH6aymZQYXIfnlqaZF9kEfeFQPmUoo2dwWtqgUvuX6ImvO0/KUdUEgMvgOke4l2o5
7GdcEFQX9r8U5UwrUn+9qQ5zlzDcyaToNrFz5UcmYyd3VhuIjM5wFP43j5X5dqMJ8CXtX6RHFEJJ
eFfJytZyJWBGm/YnrRAXNX2qVWqEdNxh8B7sKoE67ynwjwFXu/gi2q61Oi/aWXKXMR+Eww+FXLrh
f/nERkGPyVcfrBlL/GcDHJ+2gliHm9962JxkeodwNSGHLAnQ8JuAMgwulkBuIi82q2OHB3INUgwR
SbijkRfjlNP50faa7mKj02l9OScNVA7FCMW8aF2cQUsZl/StrgsY+1GcmOmaTw14LcZEyE9Uem0X
Dgkj7DoOLmgadfHPYn3xS4yhkcNcsehjoX5eTh3aurukEkJPwdqwKMkosB5cokkMsKuhptnMAV+S
3313m0rQLKRja4FBmsSJBiLV1FtoX17G+yqhWtHt3RhuQ98ISvjnjZjyUF1eAc5JhZwqAANvseLq
XZMM0glbx7m45ngqzF5qh5RCMitJkeF/xb0HKoQIk4PgBf6HZmCSNebn5c2iZ5cbfnOT10K/yX25
1f5Ml6PNiUMj7YCjALYdePQBaLFNyg13LQRVDh20Rw2fd3XtGD93PXQCvne07CEtEDBJXv1BR9ci
mK2t28hkT6amtTTM/mZQxc5C79dY4qu26os0kiQkcjcOsh8/LKMGRkW2WAjDdKvGsz69i7EQBMP4
ngmRq4OAY7TKyQj/L6lg85RaYBxDRApAE4nDcDjjSpDsELZEkpotVjc+bDKJ0R/GbKUjvhSs80xI
NW6XZuUsd/Gw6fGEqy0EZ8qhHSmNK8wi3WiKLH4JU7MJu41IxPACodGjE9SkaMZDA05K/l5d4ToY
avHgyeYkwjVBXOOrU8R3hTiG8wN7TwVlyWIEmeKU881RUI5EENobxfTRe71gwxXni1B6XH0ABbq9
l+wkkQXoJxqWw5x1FtjejG8Sd/OuE69PDIcmbVICU/77mGk++4whmZhimCXFYVWte1Db1Pe/a8iv
rnPgBcq7/LCtNJNlyGISA+yM/pWaqZbWuvEP+IHesbUMSyKiVGFbgKAJbtGwumiRdIEyCHTlW6Oo
P4cSXQm+o1VUyQzP3+UwObwFyWNmf6UmpOoHfI8fFaKKtljIW5v/Lx6XUmlArrOi23u2+/MslR8e
Y4N2MrtsTnW6WXTpWG28BecUYW35+jQi65e6BoiblHUSI0d+sazcnxr/wRC7rr971AepAZKhPHO/
TywhH61b04nptYfm8P3egCn8NaVpFpKVtNT2p5p65VXnsSSrb3990d2e+NfN1BH2NTqfYV3O53Jq
aQ6602qC/kSX9BmcHBTJOO1QdBHU4BG1WqJgKnplvjFiBDYpVpuDUSENuf52OqsCAiK9miN4F46q
m4S3s868enFFhq2UW2mrKIPyt2AY7lL3/KcFOL1v+9Ere/9j+4JQV9UMqg37PGFU3DWrTgF6GPzF
Y2hRPAJwwZf2BPoGR3paGCp71atmwyPiK0CkVR/qxs5xLLRwEQndRz2LtspI7jR/Y0oZiwWJ8lUr
uKORqpPQ6wYaFiarxPtfbxVIQe83cc+hhr1zd+CWHZkzfndKbACILXy575PMG23afr5KRbGj+QC/
sAO4hV7ldRxcDzI2l/ZrIyCas8K3WSTdBfBxQO+x+pe9H7bOjuuxurucuUUO2D5AHRj3HX+pCdLY
8zOpGj50FCTw0l5PkVHH33RmrlbP/ZPiI+1wUpB3iZxxgTZGsjQHepnEt3E9CHumkDXAI2Qd9dVT
c3Pxd4CfAQrnsdQD1Bfu5TLN4a5ZD3iPeB3YnWCQSkZCSKsSxPdCTWi994qCxeKUXcMB+5INJmX8
YjtjLFnlmzyx+l9m5iAOYqwcJGysWy1bO4hBUEl17wBrfYWPS2EdrjZUTJ4sfiwunxf04bYxK3U5
tEyjAUDftL5keuSWGnEZNIbKrSpw3h7OUV+ns0JVu0j6h5CSIC3yOnFIawv/PY+fuULd8M7mjNZQ
AO7V5fjboXWsPA96YNzw+esiLAvas6teGwSdx1yy+ohjwdQWv72Lj9PUKYRbpPYPY2BFNihvibTP
4u1SjYMxCE9wui7Ok+TQw7nxmVwOK2fyc6nvJ/TRExVEsXNObhazdC8kAAcnltR5Js7dmKYkoLkW
cmp+rHDguykVXzcPVIuLWudm9idQEfSGAAJxvJyWfIhX6UbgCzrGm+2G/w71vyNhV9oY4PaJdMRh
bhaodju64lxgy9HB0jg/9G3lzecWjvN/+cZEfeOg9omP57Xlx53FZbGXCib4KRMREPqRbzg/Tr8E
7e1R/rd2JZcp7nXn39iiQSuT3thbP8JsG3ydcobq0MpOXUX2mdyclZp9IxuOMpTKaccY6tTr6whU
qJHpcfTC/11A9xypLwzOBA0DR58ZY1t88OfSjaBmSxKaeJH8LAOjySXDcJFIzxmrtUCN56ehtVD9
EJMJzfuAPtJA0Y/nfRzJ93o4Fmoj2R55g5YD9zN/x96ujQ0ww+8a0Y7oEW2uDbnAcAavW6dFSVA0
ANrvyMdbvRVHBfLHhBa5qPYShwxwNlhut/iMKr1J6ZlpPOF0IkKT5PPkJZ1iGNqC33LpCtfVpMGH
67yheuDeq2jKHwRJpjxhjsx7Q71/O5SySDSo/B1233EhrBpCfp33waMstrIfzwVtw3PElRQxS7Gy
oWFg1NfBmWvljLK2UdyEe3PH882iHE/HgJs1qvuUMbMnvHl///gtkrjTkJ0xUVSShqAYb6y6z2xC
Tehn7PSkCP7/QgKpcYY9PjEpkezYrXQCoMN30rCGlx8ENCBIl7pwR/GkS3pPbcVm3pYLMUoSqout
oxa/RbVUcFueLHb6WQNVQ8MCsJ4i3zrahUXi+L6wIIc8n5kzNMSyp7m5O43OrA8PiL8P9JiL2X6G
UwrKCnQ1Gv0BGZ3U2vpHOsk/LkLhRoWS83BhMceNAnDMe9S37qpDWg4VZX5JXMlDy1e/FH30y3Zk
Wzma/U40V240DpJkjhz1wadx0bV7wfxnwdt3fZ9pfyNVVB2ZE0Fl/ip4Ir/myiR1OBat+SXcKRjU
5Lw9i0+vdSX7iTiz3ttU6atS8UOUeO162W5GzYeE1SKldvrlVoFAH3yslvMKLbSsKBg5NR8fkE5+
06QlxDTXxuXd7jiqga0Cz9YmRk/+esmUQFF/4hAiPD/i0tgEQDu/8GH3UYXDUSnqcouh8ixfQLcU
SB/QWfA0ddTby3/rKsRELmiwNrn6vSxW1a97Rq8tA8C6oHFdqu75+hdPCeYccNtywDScE81o9y4y
XwGV7PHGRS/x73jMUOEqniAwuhiZThlSeOZRFtT0Wy/whCDY1Gj+OdEfKbh3J0fOs1fiOY1l3tcY
+uLKx7iGmG1AZKipNPbFqNILtNzFbZFyRn5QCGC0i7dDGhH2Evs14c9/sUSzhzT6QmfZEbGISwqz
5fdEifAKE2JYbYl8KplZEwbM4lexWKpD0BVlcm4jwPtkNm8k5tCiVwxqgtm2Ikk/7CPDPStNt+mb
n7M2HI5a3jTRQ2B+Oi3C5ko+q4l7Rqacm8I4Csuyp8NpS8ciHXNgs4IGMDS1lXsuNzLHP0eDQGh9
yVYIaTQFYuDxJScE5MDROUaeKva4Y6tdr5bB4cnZyGrtj/8RRC0mjFhPm1eLoGTkqeLNSHd+++cO
UB+U9gjcqMR0ODdcmpCgeRhT8QhKAEfMeCSpughiwVDa3okHwOFPsDP4ora2NNiAcda72fZhWSlI
o0/hg9qlHJZIRMUdT7NBLsu/Vuk0tWs4UBHjc67X0kZBrCatFGvxala3Hiqu61XWFK/HRi+hIaYb
03KuYfwMkCJvU4v6IYmMBkqFGJy0/MunFYuvRbdmq6Bn7yqci+H6wk5q5W1Y2UE6yxFHe4OPsQPQ
VtPr8sh8nbsqyekwSwHiCZdJmyhlLsNcp5Ytb6V7kpKazJh4jtC5P7W9E0TOmf77idFQI6SfBHrd
TPW6aY3SxpGY6VF0F4Z5ctWil6J5BFLLxhd2ULIQBakgA1y2Q81FvQIOJP7kSUzxQZm4XwbqMfwi
MBlV3FpBuSngYbjHO0KHkX7peh1Vy0uIJqNv8bOo7v1KagN1zMiz1CgR6lNoKDRTiyETBngd9CPO
XowMHQA1KHcFHLN/NG2GqSFhiKOC50xTL02oXr73mRWAdZPVnQXtyhhgDYZXnXfMPSyFyaGzYxPB
hIVbyrlpKuxFTThiaYPShFjMRJ73oA6+GNBM4x/M21rToPi7KXs0cdG3Ekx+8I1suAW6PU62mw9I
9L9OBsqhZD7TPNBEfOGBI/5oX8XUSXKjDLFe95QRLP9BMLKc6QuR6ZBtzXQQxD+Bo0eoQsl4Yprr
n0gxw7UA5VC5BoZA6BeSvWmwLvdbrDBPepFsEuaLy3STTXOuI1LXb2bj6Alu3eAcb9/X+LDjsTDP
nu3zAJbHV1kfh4DVGs3MexRXKqmagF9a/67228z6Y7atRCUycN2RfP2iJfoGd0fX8zuMuZG6+HjJ
srmhIANJkH4rFnapWn4RGLcqUiIMBWV1MIeH/zGLN3COaLDTbO2oHl8JiW6O+uAftDhsnUs3kdDs
Yk0HpMXHu9xfq6LU+9ibA6BbIGRwmznl5taHt0qiQOq+tCU+lWwZjsrugyKLAxlvOd6ojW7/xbkD
NLSzR9mwant/qyhCn3MfG5TeErjFQPBCIGqizH4LbDYJ1LEBe2xiggdTCLRZSz/oMVbteIdftdCN
azim0mWcPR+9zn0GO332UEvKJhneRX5DXBJBB2AocMS6ezOE9RfMG0pLF5rizD8cxzebchq5j7Q6
tvQeoGdZvx84xuO+lZDvYczHvgLQ/BfxXNeLFMiwztLUNYenRUN0lz5z15LWsrxMh9dvA4D8Zf/j
8c1SHwItlmqcucCf6mClW+K940CrfN6ulyD2D+lJ+TrfhLKIuZc+48lMEyzEnx37q+zk8TNt2Mpc
H0x+qCX1WAeatk4jKQO8QCmkNpe1hbaEjCQJW3iQS+d+ukHbaexBVjf7luXDirjk2Xu2sFpOs/CG
dHwuJYA8j4dJXuerMH1zIk8c9jScIwuI714FQHA6AJLXEoXbBtt1tr+XNd52NLCK/xrzpjDfuZOU
RwmhFOzCzGQN9p3S834Pg3ELaCBO/ftp1eYwEiyhCAiAoN7fDB0Gf4+XoLhPAdpvToo9cqfYPWDh
4T0WfmPxAknx4xL9EN/HQYNhFXx93F0XHJRSjfQPj6ozLA9E4fQ+e86Ho1j7WuUWNACpJlWGtAqU
BaSwxNae0Gr+OrCecp94Y9uUXZgnI7wxku23rqPbY16Q68b5p+RZRDR6nZdGoNfLs8/bEQ6dGxDG
2eCnr4bI8fFprxYouKrzHmhGfbBpF7WmVepjLwInSdi/Tryn+hnqevFE/6+lywpc/QOCSHRNTLHO
YZ4PgMAZsdHL3aefEdD8M+oh1FHhysS6CbYDK53xyKDxWSgQbvDFBG4rwOv2yDj7JjK37437tK/4
e5OEfbgsfuNuGSu26eCjRJ6IXzl7TiUKyloIDPgnjGL2UHB2Y9iDTRUXEfBVxNgW62VY3eSlFmTY
bzSg4y3mQczgMPJr3946wlFDrJGkMz8u74Yh/njt3DpWC5ySMvLcMDN11orXKyB0yWwZsKPA6q2A
3f2H+toMGRFzBwnZejv0F/6vekSkqvozLPu13sQ7A/9wo3iw2g+7/05hmgyJH8scioYvSZRMjbJd
JJcXQv1L/83UHjH7Mq7nYq+tC7dhtvgbB9E9wLkaiyVE8vF/wTuOxg3mPsnpg/wIGKoruo992xFX
bPekRVoIb9+gZ2eO1+ES4OtzFRt2ibiXxtWnTvyNS60em9US+KDcC+5GKNG/I93Y1G/CpmW7Bnxk
tzisN4lkZXacqFlegxJ/MpUbchVXRc2GlFGpFcXCIeXL2XjseC09V5RS3pCl+26FsEO9tfglD0dU
AGRXztUy1ZQdm7MKPu2lzpI4CclWCOm18WhnF+Jr4kAWGHZfCP74rLT2/DoT4YT96e5joi2lVgaS
IDad4F/tBJKWOmpEu6JKV9FdjDEc9CqF5DJt3vQ6UrgOlxtpm41GQmIJrqnPlN0y83VXuMJ+eCzj
XuydXX5OeX0SGhpd+rNwt0DL9EIWNF9OUpAE4DUL1pitmy0iIkQPLXCt5eXqYeCSRjkixLPQBYdF
DyYgMi1YK989IFNHosE9Vswm3/N3dCoeBfsFqG1CYHXktoh/ZbJ57U7Yf+dS6RHReoQs44G1laIq
wOrsPR47KVuvizKCui8F8iaLORqR+XcPUJHbgJLZ1PLUOY6TWYmvpacN3BIfkNSPyX1VeCirc6B4
y1Mcz4WFs6e9YYDWG8RwlpNSIONKnOxX2x9oLfY=
`protect end_protected
